// controller.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module controller (
		input  wire        adc2_i2c_scl_in,                                          //     adc2_i2c.scl_in
		input  wire        adc2_i2c_sda_in,                                          //             .sda_in
		output wire        adc2_i2c_scl_oe,                                          //             .scl_oe
		output wire        adc2_i2c_sda_oe,                                          //             .sda_oe
		input  wire        clk_100mhz_clk,                                           //   clk_100mhz.clk
		input  wire        clk_sys_clk,                                              //      clk_sys.clk
		input  wire        host_spi_mosi_to_the_spislave_inst_for_spichain,          //     host_spi.mosi_to_the_spislave_inst_for_spichain
		input  wire        host_spi_nss_to_the_spislave_inst_for_spichain,           //             .nss_to_the_spislave_inst_for_spichain
		inout  wire        host_spi_miso_to_and_from_the_spislave_inst_for_spichain, //             .miso_to_and_from_the_spislave_inst_for_spichain
		input  wire        host_spi_sclk_to_the_spislave_inst_for_spichain,          //             .sclk_to_the_spislave_inst_for_spichain
		output wire        imu_spi_mosi,                                             //      imu_spi.mosi
		input  wire        imu_spi_miso,                                             //             .miso
		output wire        imu_spi_sclk,                                             //             .sclk
		output wire        imu_spi_cs_n,                                             //             .cs_n
		input  wire        imu_spi_int_n,                                            //             .int_n
		output wire        mc5_fault_fault,                                          //    mc5_fault.fault
		output wire        mc5_fault_brake,                                          //             .brake
		output wire [15:0] mc5_pwm_data,                                             //      mc5_pwm.data
		output wire        mc5_pwm_valid,                                            //             .valid
		input  wire        mc5_pwm_ready,                                            //             .ready
		input  wire        mc5_status_driver_otw_n,                                  //   mc5_status.driver_otw_n
		input  wire        mc5_status_driver_fault_n,                                //             .driver_fault_n
		input  wire        mc5_status_hall_fault_n,                                  //             .hall_fault_n
		input  wire        pio_0_export,                                             //        pio_0.export
		input  wire [31:0] pio_1_export,                                             //        pio_1.export
		output wire [9:0]  pio_2_export,                                             //        pio_2.export
		input  wire        reset_100mhz_reset_n,                                     // reset_100mhz.reset_n
		input  wire        reset_ext_reset,                                          //    reset_ext.reset
		input  wire        reset_sys_reset_n,                                        //    reset_sys.reset_n
		output wire        uart_txd,                                                 //         uart.txd
		input  wire [15:0] vc_encoder_encoder_1_data,                                //   vc_encoder.encoder_1_data
		input  wire [15:0] vc_encoder_encoder_2_data,                                //             .encoder_2_data
		input  wire [15:0] vc_encoder_encoder_3_data,                                //             .encoder_3_data
		input  wire [15:0] vc_encoder_encoder_4_data,                                //             .encoder_4_data
		output wire        vc_fault_fault,                                           //     vc_fault.fault
		output wire [3:0]  vc_fault_brake,                                           //             .brake
		input  wire [31:0] vc_imeas1_data,                                           //    vc_imeas1.data
		input  wire        vc_imeas1_valid,                                          //             .valid
		input  wire [31:0] vc_imeas2_data,                                           //    vc_imeas2.data
		input  wire        vc_imeas2_valid,                                          //             .valid
		input  wire [31:0] vc_imeas3_data,                                           //    vc_imeas3.data
		input  wire        vc_imeas3_valid,                                          //             .valid
		input  wire [31:0] vc_imeas4_data,                                           //    vc_imeas4.data
		input  wire        vc_imeas4_valid,                                          //             .valid
		output wire [31:0] vc_iref1_data,                                            //     vc_iref1.data
		output wire        vc_iref1_valid,                                           //             .valid
		output wire [31:0] vc_iref2_data,                                            //     vc_iref2.data
		output wire        vc_iref2_valid,                                           //             .valid
		output wire [31:0] vc_iref3_data,                                            //     vc_iref3.data
		output wire        vc_iref3_valid,                                           //             .valid
		output wire [31:0] vc_iref4_data,                                            //     vc_iref4.data
		output wire        vc_iref4_valid,                                           //             .valid
		output wire [15:0] vc_param_kp,                                              //     vc_param.kp
		output wire [15:0] vc_param_ki,                                              //             .ki
		input  wire [3:0]  vc_status_driver_otw_n,                                   //    vc_status.driver_otw_n
		input  wire [3:0]  vc_status_driver_fault_n,                                 //             .driver_fault_n
		input  wire [3:0]  vc_status_hall_fault_n,                                   //             .hall_fault_n
		input  wire [3:0]  vc_status_encoder_fault_n,                                //             .encoder_fault_n
		input  wire [3:0]  vc_status_pos_error,                                      //             .pos_error
		input  wire [3:0]  vc_status_pos_uncertain                                   //             .pos_uncertain
	);

	wire          vic_0_interrupt_controller_out_valid;                                         // vic_0:interrupt_controller_out_valid -> nios_0:eic_port_valid
	wire   [44:0] vic_0_interrupt_controller_out_data;                                          // vic_0:interrupt_controller_out_data -> nios_0:eic_port_data
	wire          dc_fifo_0_out_valid;                                                          // dc_fifo_0:out_valid -> avalon_st_uart_tx_0:sink_valid
	wire    [7:0] dc_fifo_0_out_data;                                                           // dc_fifo_0:out_data -> avalon_st_uart_tx_0:sink_data
	wire          dc_fifo_0_out_ready;                                                          // avalon_st_uart_tx_0:sink_ready -> dc_fifo_0:out_ready
	wire          st_packets_to_bytes_0_out_bytes_stream_valid;                                 // st_packets_to_bytes_0:out_valid -> dc_fifo_0:in_valid
	wire    [7:0] st_packets_to_bytes_0_out_bytes_stream_data;                                  // st_packets_to_bytes_0:out_data -> dc_fifo_0:in_data
	wire          st_packets_to_bytes_0_out_bytes_stream_ready;                                 // dc_fifo_0:in_ready -> st_packets_to_bytes_0:out_ready
	wire          msgdma_0_st_source_valid;                                                     // msgdma_0:st_source_valid -> st_packets_to_bytes_0:in_valid
	wire    [7:0] msgdma_0_st_source_data;                                                      // msgdma_0:st_source_data -> st_packets_to_bytes_0:in_data
	wire          msgdma_0_st_source_ready;                                                     // st_packets_to_bytes_0:in_ready -> msgdma_0:st_source_ready
	wire    [7:0] msgdma_0_st_source_channel;                                                   // msgdma_0:st_source_channel -> st_packets_to_bytes_0:in_channel
	wire          msgdma_0_st_source_startofpacket;                                             // msgdma_0:st_source_startofpacket -> st_packets_to_bytes_0:in_startofpacket
	wire          msgdma_0_st_source_endofpacket;                                               // msgdma_0:st_source_endofpacket -> st_packets_to_bytes_0:in_endofpacket
	wire          spim_0_external_sclk;                                                         // spim_0:SCLK -> imu_spim:SCLK
	wire          spim_0_external_ss_n;                                                         // spim_0:SS_n -> imu_spim:SS_n
	wire          imu_spim_spis_miso;                                                           // imu_spim:MISO -> spim_0:MISO
	wire          spim_0_external_mosi;                                                         // spim_0:MOSI -> imu_spim:MOSI
	wire          nios_0_custom_instruction_master_readra;                                      // nios_0:E_ci_combo_readra -> nios_0_custom_instruction_master_translator:ci_slave_readra
	wire          nios_0_custom_instruction_master_readrb;                                      // nios_0:E_ci_combo_readrb -> nios_0_custom_instruction_master_translator:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_multi_b;                                     // nios_0:A_ci_multi_b -> nios_0_custom_instruction_master_translator:ci_slave_multi_b
	wire    [4:0] nios_0_custom_instruction_master_multi_c;                                     // nios_0:A_ci_multi_c -> nios_0_custom_instruction_master_translator:ci_slave_multi_c
	wire          nios_0_custom_instruction_master_reset_req;                                   // nios_0:A_ci_multi_reset_req -> nios_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire    [4:0] nios_0_custom_instruction_master_multi_a;                                     // nios_0:A_ci_multi_a -> nios_0_custom_instruction_master_translator:ci_slave_multi_a
	wire   [31:0] nios_0_custom_instruction_master_result;                                      // nios_0_custom_instruction_master_translator:ci_slave_result -> nios_0:E_ci_combo_result
	wire   [31:0] nios_0_custom_instruction_master_datab;                                       // nios_0:E_ci_combo_datab -> nios_0_custom_instruction_master_translator:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_dataa;                                       // nios_0:E_ci_combo_dataa -> nios_0_custom_instruction_master_translator:ci_slave_dataa
	wire          nios_0_custom_instruction_master_writerc;                                     // nios_0:E_ci_combo_writerc -> nios_0_custom_instruction_master_translator:ci_slave_writerc
	wire   [31:0] nios_0_custom_instruction_master_multi_dataa;                                 // nios_0:A_ci_multi_dataa -> nios_0_custom_instruction_master_translator:ci_slave_multi_dataa
	wire          nios_0_custom_instruction_master_multi_writerc;                               // nios_0:A_ci_multi_writerc -> nios_0_custom_instruction_master_translator:ci_slave_multi_writerc
	wire    [4:0] nios_0_custom_instruction_master_a;                                           // nios_0:E_ci_combo_a -> nios_0_custom_instruction_master_translator:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_b;                                           // nios_0:E_ci_combo_b -> nios_0_custom_instruction_master_translator:ci_slave_b
	wire   [31:0] nios_0_custom_instruction_master_multi_result;                                // nios_0_custom_instruction_master_translator:ci_slave_multi_result -> nios_0:A_ci_multi_result
	wire          nios_0_custom_instruction_master_clk;                                         // nios_0:A_ci_multi_clock -> nios_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire   [31:0] nios_0_custom_instruction_master_multi_datab;                                 // nios_0:A_ci_multi_datab -> nios_0_custom_instruction_master_translator:ci_slave_multi_datab
	wire    [4:0] nios_0_custom_instruction_master_c;                                           // nios_0:E_ci_combo_c -> nios_0_custom_instruction_master_translator:ci_slave_c
	wire   [31:0] nios_0_custom_instruction_master_ipending;                                    // nios_0:E_ci_combo_ipending -> nios_0_custom_instruction_master_translator:ci_slave_ipending
	wire          nios_0_custom_instruction_master_start;                                       // nios_0:A_ci_multi_start -> nios_0_custom_instruction_master_translator:ci_slave_multi_start
	wire          nios_0_custom_instruction_master_done;                                        // nios_0_custom_instruction_master_translator:ci_slave_multi_done -> nios_0:A_ci_multi_done
	wire    [7:0] nios_0_custom_instruction_master_n;                                           // nios_0:E_ci_combo_n -> nios_0_custom_instruction_master_translator:ci_slave_n
	wire          nios_0_custom_instruction_master_estatus;                                     // nios_0:E_ci_combo_estatus -> nios_0_custom_instruction_master_translator:ci_slave_estatus
	wire          nios_0_custom_instruction_master_clk_en;                                      // nios_0:A_ci_multi_clk_en -> nios_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire          nios_0_custom_instruction_master_reset;                                       // nios_0:A_ci_multi_reset -> nios_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire          nios_0_custom_instruction_master_multi_readrb;                                // nios_0:A_ci_multi_readrb -> nios_0_custom_instruction_master_translator:ci_slave_multi_readrb
	wire          nios_0_custom_instruction_master_multi_readra;                                // nios_0:A_ci_multi_readra -> nios_0_custom_instruction_master_translator:ci_slave_multi_readra
	wire    [7:0] nios_0_custom_instruction_master_multi_n;                                     // nios_0:A_ci_multi_n -> nios_0_custom_instruction_master_translator:ci_slave_multi_n
	wire   [31:0] nios_0_custom_instruction_master_translator_comb_ci_master_result;            // nios_0_custom_instruction_master_comb_xconnect:ci_slave_result -> nios_0_custom_instruction_master_translator:comb_ci_master_result
	wire          nios_0_custom_instruction_master_translator_comb_ci_master_readra;            // nios_0_custom_instruction_master_translator:comb_ci_master_readra -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire    [4:0] nios_0_custom_instruction_master_translator_comb_ci_master_a;                 // nios_0_custom_instruction_master_translator:comb_ci_master_a -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_translator_comb_ci_master_b;                 // nios_0_custom_instruction_master_translator:comb_ci_master_b -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_b
	wire          nios_0_custom_instruction_master_translator_comb_ci_master_readrb;            // nios_0_custom_instruction_master_translator:comb_ci_master_readrb -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_translator_comb_ci_master_c;                 // nios_0_custom_instruction_master_translator:comb_ci_master_c -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_c
	wire          nios_0_custom_instruction_master_translator_comb_ci_master_estatus;           // nios_0_custom_instruction_master_translator:comb_ci_master_estatus -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire   [31:0] nios_0_custom_instruction_master_translator_comb_ci_master_ipending;          // nios_0_custom_instruction_master_translator:comb_ci_master_ipending -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire   [31:0] nios_0_custom_instruction_master_translator_comb_ci_master_datab;             // nios_0_custom_instruction_master_translator:comb_ci_master_datab -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_translator_comb_ci_master_dataa;             // nios_0_custom_instruction_master_translator:comb_ci_master_dataa -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire          nios_0_custom_instruction_master_translator_comb_ci_master_writerc;           // nios_0_custom_instruction_master_translator:comb_ci_master_writerc -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire    [7:0] nios_0_custom_instruction_master_translator_comb_ci_master_n;                 // nios_0_custom_instruction_master_translator:comb_ci_master_n -> nios_0_custom_instruction_master_comb_xconnect:ci_slave_n
	wire   [31:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_result;             // nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios_0_custom_instruction_master_comb_xconnect:ci_master0_result
	wire          nios_0_custom_instruction_master_comb_xconnect_ci_master0_readra;             // nios_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire    [4:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_a;                  // nios_0_custom_instruction_master_comb_xconnect:ci_master0_a -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_b;                  // nios_0_custom_instruction_master_comb_xconnect:ci_master0_b -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire          nios_0_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // nios_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_c;                  // nios_0_custom_instruction_master_comb_xconnect:ci_master0_c -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire          nios_0_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // nios_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire   [31:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // nios_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire   [31:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_datab;              // nios_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // nios_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire          nios_0_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // nios_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire    [7:0] nios_0_custom_instruction_master_comb_xconnect_ci_master0_n;                  // nios_0_custom_instruction_master_comb_xconnect:ci_master0_n -> nios_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire   [31:0] nios_0_custom_instruction_master_comb_slave_translator0_ci_master_result;     // fpu_0:s1_result -> nios_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire   [31:0] nios_0_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // nios_0_custom_instruction_master_comb_slave_translator0:ci_master_datab -> fpu_0:s1_datab
	wire   [31:0] nios_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // nios_0_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> fpu_0:s1_dataa
	wire    [3:0] nios_0_custom_instruction_master_comb_slave_translator0_ci_master_n;          // nios_0_custom_instruction_master_comb_slave_translator0:ci_master_n -> fpu_0:s1_n
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_readra;           // nios_0_custom_instruction_master_translator:multi_ci_master_readra -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire    [4:0] nios_0_custom_instruction_master_translator_multi_ci_master_a;                // nios_0_custom_instruction_master_translator:multi_ci_master_a -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_translator_multi_ci_master_b;                // nios_0_custom_instruction_master_translator:multi_ci_master_b -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_clk;              // nios_0_custom_instruction_master_translator:multi_ci_master_clk -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_readrb;           // nios_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_translator_multi_ci_master_c;                // nios_0_custom_instruction_master_translator:multi_ci_master_c -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_start;            // nios_0_custom_instruction_master_translator:multi_ci_master_start -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_reset_req;        // nios_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_done;             // nios_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios_0_custom_instruction_master_translator:multi_ci_master_done
	wire    [7:0] nios_0_custom_instruction_master_translator_multi_ci_master_n;                // nios_0_custom_instruction_master_translator:multi_ci_master_n -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire   [31:0] nios_0_custom_instruction_master_translator_multi_ci_master_result;           // nios_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios_0_custom_instruction_master_translator:multi_ci_master_result
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_clk_en;           // nios_0_custom_instruction_master_translator:multi_ci_master_clken -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire   [31:0] nios_0_custom_instruction_master_translator_multi_ci_master_datab;            // nios_0_custom_instruction_master_translator:multi_ci_master_datab -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_translator_multi_ci_master_dataa;            // nios_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_reset;            // nios_0_custom_instruction_master_translator:multi_ci_master_reset -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire          nios_0_custom_instruction_master_translator_multi_ci_master_writerc;          // nios_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_readra;            // nios_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_a;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_b;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // nios_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_c;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk;               // nios_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // nios_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_start;             // nios_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // nios_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_done;              // nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire    [7:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_n;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_result;            // nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // nios_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // nios_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_datab;             // nios_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // nios_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset;             // nios_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // nios_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire   [31:0] nios_0_custom_instruction_master_multi_slave_translator0_ci_master_result;    // float32to16_0:slave_result -> nios_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire          nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // nios_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> float32to16_0:slave_clk
	wire          nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // nios_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> float32to16_0:slave_clk_en
	wire   [31:0] nios_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // nios_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> float32to16_0:slave_dataa
	wire          nios_0_custom_instruction_master_multi_slave_translator0_ci_master_start;     // nios_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> float32to16_0:slave_start
	wire          nios_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // nios_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> float32to16_0:slave_reset
	wire          nios_0_custom_instruction_master_multi_slave_translator0_ci_master_done;      // float32to16_0:slave_done -> nios_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_readra;            // nios_0_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_a;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master1_a -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_b;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master1_b -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_readrb;            // nios_0_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire    [4:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_c;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master1_c -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk;               // nios_0_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_ipending;          // nios_0_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_start;             // nios_0_custom_instruction_master_multi_xconnect:ci_master1_start -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req;         // nios_0_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_done;              // nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios_0_custom_instruction_master_multi_xconnect:ci_master1_done
	wire    [7:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_n;                 // nios_0_custom_instruction_master_multi_xconnect:ci_master1_n -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_result;            // nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios_0_custom_instruction_master_multi_xconnect:ci_master1_result
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_estatus;           // nios_0_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en;            // nios_0_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_datab;             // nios_0_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire   [31:0] nios_0_custom_instruction_master_multi_xconnect_ci_master1_dataa;             // nios_0_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset;             // nios_0_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire          nios_0_custom_instruction_master_multi_xconnect_ci_master1_writerc;           // nios_0_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios_0_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire   [31:0] nios_0_custom_instruction_master_multi_slave_translator1_ci_master_result;    // fpu_0:s2_result -> nios_0_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk;       // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_clk -> fpu_0:s2_clk
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en;    // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_clken -> fpu_0:s2_clk_en
	wire   [31:0] nios_0_custom_instruction_master_multi_slave_translator1_ci_master_datab;     // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_datab -> fpu_0:s2_datab
	wire   [31:0] nios_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa;     // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> fpu_0:s2_dataa
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_start;     // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_start -> fpu_0:s2_start
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset;     // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_reset -> fpu_0:s2_reset
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset_req; // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_reset_req -> fpu_0:s2_reset_req
	wire          nios_0_custom_instruction_master_multi_slave_translator1_ci_master_done;      // fpu_0:s2_done -> nios_0_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire    [2:0] nios_0_custom_instruction_master_multi_slave_translator1_ci_master_n;         // nios_0_custom_instruction_master_multi_slave_translator1:ci_master_n -> fpu_0:s2_n
	wire   [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata;                // mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata -> spi_slave_to_avalon_mm_master_bridge_0:readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire          spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest;             // mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest -> spi_slave_to_avalon_mm_master_bridge_0:waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire   [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address;                 // spi_slave_to_avalon_mm_master_bridge_0:address_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address
	wire    [3:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable;              // spi_slave_to_avalon_mm_master_bridge_0:byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable
	wire          spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read;                    // spi_slave_to_avalon_mm_master_bridge_0:read_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read
	wire          spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid;           // mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid -> spi_slave_to_avalon_mm_master_bridge_0:readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire          spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write;                   // spi_slave_to_avalon_mm_master_bridge_0:write_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write
	wire   [31:0] spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata;               // spi_slave_to_avalon_mm_master_bridge_0:writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata
	wire   [31:0] mm_interconnect_0_mm_bridge_2_s0_readdata;                                    // mm_bridge_2:s0_readdata -> mm_interconnect_0:mm_bridge_2_s0_readdata
	wire          mm_interconnect_0_mm_bridge_2_s0_waitrequest;                                 // mm_bridge_2:s0_waitrequest -> mm_interconnect_0:mm_bridge_2_s0_waitrequest
	wire          mm_interconnect_0_mm_bridge_2_s0_debugaccess;                                 // mm_interconnect_0:mm_bridge_2_s0_debugaccess -> mm_bridge_2:s0_debugaccess
	wire   [14:0] mm_interconnect_0_mm_bridge_2_s0_address;                                     // mm_interconnect_0:mm_bridge_2_s0_address -> mm_bridge_2:s0_address
	wire          mm_interconnect_0_mm_bridge_2_s0_read;                                        // mm_interconnect_0:mm_bridge_2_s0_read -> mm_bridge_2:s0_read
	wire    [3:0] mm_interconnect_0_mm_bridge_2_s0_byteenable;                                  // mm_interconnect_0:mm_bridge_2_s0_byteenable -> mm_bridge_2:s0_byteenable
	wire          mm_interconnect_0_mm_bridge_2_s0_readdatavalid;                               // mm_bridge_2:s0_readdatavalid -> mm_interconnect_0:mm_bridge_2_s0_readdatavalid
	wire          mm_interconnect_0_mm_bridge_2_s0_write;                                       // mm_interconnect_0:mm_bridge_2_s0_write -> mm_bridge_2:s0_write
	wire   [31:0] mm_interconnect_0_mm_bridge_2_s0_writedata;                                   // mm_interconnect_0:mm_bridge_2_s0_writedata -> mm_bridge_2:s0_writedata
	wire    [0:0] mm_interconnect_0_mm_bridge_2_s0_burstcount;                                  // mm_interconnect_0:mm_bridge_2_s0_burstcount -> mm_bridge_2:s0_burstcount
	wire          mm_interconnect_0_data_ram_1_s2_chipselect;                                   // mm_interconnect_0:data_ram_1_s2_chipselect -> data_ram_1:chipselect2
	wire   [31:0] mm_interconnect_0_data_ram_1_s2_readdata;                                     // data_ram_1:readdata2 -> mm_interconnect_0:data_ram_1_s2_readdata
	wire    [7:0] mm_interconnect_0_data_ram_1_s2_address;                                      // mm_interconnect_0:data_ram_1_s2_address -> data_ram_1:address2
	wire    [3:0] mm_interconnect_0_data_ram_1_s2_byteenable;                                   // mm_interconnect_0:data_ram_1_s2_byteenable -> data_ram_1:byteenable2
	wire          mm_interconnect_0_data_ram_1_s2_write;                                        // mm_interconnect_0:data_ram_1_s2_write -> data_ram_1:write2
	wire   [31:0] mm_interconnect_0_data_ram_1_s2_writedata;                                    // mm_interconnect_0:data_ram_1_s2_writedata -> data_ram_1:writedata2
	wire          mm_interconnect_0_data_ram_1_s2_clken;                                        // mm_interconnect_0:data_ram_1_s2_clken -> data_ram_1:clken2
	wire   [31:0] nios_0_data_master_readdata;                                                  // mm_interconnect_1:nios_0_data_master_readdata -> nios_0:d_readdata
	wire          nios_0_data_master_waitrequest;                                               // mm_interconnect_1:nios_0_data_master_waitrequest -> nios_0:d_waitrequest
	wire          nios_0_data_master_debugaccess;                                               // nios_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios_0_data_master_debugaccess
	wire   [15:0] nios_0_data_master_address;                                                   // nios_0:d_address -> mm_interconnect_1:nios_0_data_master_address
	wire    [3:0] nios_0_data_master_byteenable;                                                // nios_0:d_byteenable -> mm_interconnect_1:nios_0_data_master_byteenable
	wire          nios_0_data_master_read;                                                      // nios_0:d_read -> mm_interconnect_1:nios_0_data_master_read
	wire          nios_0_data_master_write;                                                     // nios_0:d_write -> mm_interconnect_1:nios_0_data_master_write
	wire   [31:0] nios_0_data_master_writedata;                                                 // nios_0:d_writedata -> mm_interconnect_1:nios_0_data_master_writedata
	wire   [31:0] nios_0_instruction_master_readdata;                                           // mm_interconnect_1:nios_0_instruction_master_readdata -> nios_0:i_readdata
	wire          nios_0_instruction_master_waitrequest;                                        // mm_interconnect_1:nios_0_instruction_master_waitrequest -> nios_0:i_waitrequest
	wire   [15:0] nios_0_instruction_master_address;                                            // nios_0:i_address -> mm_interconnect_1:nios_0_instruction_master_address
	wire          nios_0_instruction_master_read;                                               // nios_0:i_read -> mm_interconnect_1:nios_0_instruction_master_read
	wire   [31:0] mm_interconnect_1_nios_0_debug_mem_slave_readdata;                            // nios_0:debug_mem_slave_readdata -> mm_interconnect_1:nios_0_debug_mem_slave_readdata
	wire          mm_interconnect_1_nios_0_debug_mem_slave_waitrequest;                         // nios_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_1_nios_0_debug_mem_slave_debugaccess;                         // mm_interconnect_1:nios_0_debug_mem_slave_debugaccess -> nios_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_1_nios_0_debug_mem_slave_address;                             // mm_interconnect_1:nios_0_debug_mem_slave_address -> nios_0:debug_mem_slave_address
	wire          mm_interconnect_1_nios_0_debug_mem_slave_read;                                // mm_interconnect_1:nios_0_debug_mem_slave_read -> nios_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_1_nios_0_debug_mem_slave_byteenable;                          // mm_interconnect_1:nios_0_debug_mem_slave_byteenable -> nios_0:debug_mem_slave_byteenable
	wire          mm_interconnect_1_nios_0_debug_mem_slave_write;                               // mm_interconnect_1:nios_0_debug_mem_slave_write -> nios_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_1_nios_0_debug_mem_slave_writedata;                           // mm_interconnect_1:nios_0_debug_mem_slave_writedata -> nios_0:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_1_mm_bridge_0_s0_readdata;                                    // mm_bridge_0:s0_readdata -> mm_interconnect_1:mm_bridge_0_s0_readdata
	wire          mm_interconnect_1_mm_bridge_0_s0_waitrequest;                                 // mm_bridge_0:s0_waitrequest -> mm_interconnect_1:mm_bridge_0_s0_waitrequest
	wire          mm_interconnect_1_mm_bridge_0_s0_debugaccess;                                 // mm_interconnect_1:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire   [12:0] mm_interconnect_1_mm_bridge_0_s0_address;                                     // mm_interconnect_1:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire          mm_interconnect_1_mm_bridge_0_s0_read;                                        // mm_interconnect_1:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire    [3:0] mm_interconnect_1_mm_bridge_0_s0_byteenable;                                  // mm_interconnect_1:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire          mm_interconnect_1_mm_bridge_0_s0_readdatavalid;                               // mm_bridge_0:s0_readdatavalid -> mm_interconnect_1:mm_bridge_0_s0_readdatavalid
	wire          mm_interconnect_1_mm_bridge_0_s0_write;                                       // mm_interconnect_1:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire   [31:0] mm_interconnect_1_mm_bridge_0_s0_writedata;                                   // mm_interconnect_1:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire    [0:0] mm_interconnect_1_mm_bridge_0_s0_burstcount;                                  // mm_interconnect_1:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire   [31:0] mm_interconnect_1_mm_bridge_1_s0_readdata;                                    // mm_bridge_1:s0_readdata -> mm_interconnect_1:mm_bridge_1_s0_readdata
	wire          mm_interconnect_1_mm_bridge_1_s0_waitrequest;                                 // mm_bridge_1:s0_waitrequest -> mm_interconnect_1:mm_bridge_1_s0_waitrequest
	wire          mm_interconnect_1_mm_bridge_1_s0_debugaccess;                                 // mm_interconnect_1:mm_bridge_1_s0_debugaccess -> mm_bridge_1:s0_debugaccess
	wire   [12:0] mm_interconnect_1_mm_bridge_1_s0_address;                                     // mm_interconnect_1:mm_bridge_1_s0_address -> mm_bridge_1:s0_address
	wire          mm_interconnect_1_mm_bridge_1_s0_read;                                        // mm_interconnect_1:mm_bridge_1_s0_read -> mm_bridge_1:s0_read
	wire    [3:0] mm_interconnect_1_mm_bridge_1_s0_byteenable;                                  // mm_interconnect_1:mm_bridge_1_s0_byteenable -> mm_bridge_1:s0_byteenable
	wire          mm_interconnect_1_mm_bridge_1_s0_readdatavalid;                               // mm_bridge_1:s0_readdatavalid -> mm_interconnect_1:mm_bridge_1_s0_readdatavalid
	wire          mm_interconnect_1_mm_bridge_1_s0_write;                                       // mm_interconnect_1:mm_bridge_1_s0_write -> mm_bridge_1:s0_write
	wire   [31:0] mm_interconnect_1_mm_bridge_1_s0_writedata;                                   // mm_interconnect_1:mm_bridge_1_s0_writedata -> mm_bridge_1:s0_writedata
	wire    [0:0] mm_interconnect_1_mm_bridge_1_s0_burstcount;                                  // mm_interconnect_1:mm_bridge_1_s0_burstcount -> mm_bridge_1:s0_burstcount
	wire          mm_interconnect_1_instruction_rom_0_s1_chipselect;                            // mm_interconnect_1:instruction_rom_0_s1_chipselect -> instruction_rom_0:chipselect
	wire   [31:0] mm_interconnect_1_instruction_rom_0_s1_readdata;                              // instruction_rom_0:readdata -> mm_interconnect_1:instruction_rom_0_s1_readdata
	wire   [12:0] mm_interconnect_1_instruction_rom_0_s1_address;                               // mm_interconnect_1:instruction_rom_0_s1_address -> instruction_rom_0:address
	wire    [3:0] mm_interconnect_1_instruction_rom_0_s1_byteenable;                            // mm_interconnect_1:instruction_rom_0_s1_byteenable -> instruction_rom_0:byteenable
	wire          mm_interconnect_1_instruction_rom_0_s1_write;                                 // mm_interconnect_1:instruction_rom_0_s1_write -> instruction_rom_0:write
	wire   [31:0] mm_interconnect_1_instruction_rom_0_s1_writedata;                             // mm_interconnect_1:instruction_rom_0_s1_writedata -> instruction_rom_0:writedata
	wire          mm_interconnect_1_instruction_rom_0_s1_clken;                                 // mm_interconnect_1:instruction_rom_0_s1_clken -> instruction_rom_0:clken
	wire          mm_interconnect_1_data_ram_0_s1_chipselect;                                   // mm_interconnect_1:data_ram_0_s1_chipselect -> data_ram_0:chipselect
	wire   [31:0] mm_interconnect_1_data_ram_0_s1_readdata;                                     // data_ram_0:readdata -> mm_interconnect_1:data_ram_0_s1_readdata
	wire    [9:0] mm_interconnect_1_data_ram_0_s1_address;                                      // mm_interconnect_1:data_ram_0_s1_address -> data_ram_0:address
	wire    [3:0] mm_interconnect_1_data_ram_0_s1_byteenable;                                   // mm_interconnect_1:data_ram_0_s1_byteenable -> data_ram_0:byteenable
	wire          mm_interconnect_1_data_ram_0_s1_write;                                        // mm_interconnect_1:data_ram_0_s1_write -> data_ram_0:write
	wire   [31:0] mm_interconnect_1_data_ram_0_s1_writedata;                                    // mm_interconnect_1:data_ram_0_s1_writedata -> data_ram_0:writedata
	wire          mm_interconnect_1_data_ram_0_s1_clken;                                        // mm_interconnect_1:data_ram_0_s1_clken -> data_ram_0:clken
	wire          mm_interconnect_1_data_ram_1_s1_chipselect;                                   // mm_interconnect_1:data_ram_1_s1_chipselect -> data_ram_1:chipselect
	wire   [31:0] mm_interconnect_1_data_ram_1_s1_readdata;                                     // data_ram_1:readdata -> mm_interconnect_1:data_ram_1_s1_readdata
	wire    [7:0] mm_interconnect_1_data_ram_1_s1_address;                                      // mm_interconnect_1:data_ram_1_s1_address -> data_ram_1:address
	wire    [3:0] mm_interconnect_1_data_ram_1_s1_byteenable;                                   // mm_interconnect_1:data_ram_1_s1_byteenable -> data_ram_1:byteenable
	wire          mm_interconnect_1_data_ram_1_s1_write;                                        // mm_interconnect_1:data_ram_1_s1_write -> data_ram_1:write
	wire   [31:0] mm_interconnect_1_data_ram_1_s1_writedata;                                    // mm_interconnect_1:data_ram_1_s1_writedata -> data_ram_1:writedata
	wire          mm_interconnect_1_data_ram_1_s1_clken;                                        // mm_interconnect_1:data_ram_1_s1_clken -> data_ram_1:clken
	wire          mm_bridge_0_m0_waitrequest;                                                   // mm_interconnect_2:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [31:0] mm_bridge_0_m0_readdata;                                                      // mm_interconnect_2:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                                   // mm_bridge_0:m0_debugaccess -> mm_interconnect_2:mm_bridge_0_m0_debugaccess
	wire   [12:0] mm_bridge_0_m0_address;                                                       // mm_bridge_0:m0_address -> mm_interconnect_2:mm_bridge_0_m0_address
	wire          mm_bridge_0_m0_read;                                                          // mm_bridge_0:m0_read -> mm_interconnect_2:mm_bridge_0_m0_read
	wire    [3:0] mm_bridge_0_m0_byteenable;                                                    // mm_bridge_0:m0_byteenable -> mm_interconnect_2:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                                 // mm_interconnect_2:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [31:0] mm_bridge_0_m0_writedata;                                                     // mm_bridge_0:m0_writedata -> mm_interconnect_2:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                                         // mm_bridge_0:m0_write -> mm_interconnect_2:mm_bridge_0_m0_write
	wire    [0:0] mm_bridge_0_m0_burstcount;                                                    // mm_bridge_0:m0_burstcount -> mm_interconnect_2:mm_bridge_0_m0_burstcount
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect;                   // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata;                     // jtag_uart_0:av_readdata -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest;                  // jtag_uart_0:av_waitrequest -> mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address;                      // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read;                         // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write;                        // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata;                    // mm_interconnect_2:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [31:0] mm_interconnect_2_sysid_qsys_0_control_slave_readdata;                        // sysid_qsys_0:readdata -> mm_interconnect_2:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_2_sysid_qsys_0_control_slave_address;                         // mm_interconnect_2:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_2_performance_counter_0_control_slave_readdata;               // performance_counter_0:readdata -> mm_interconnect_2:performance_counter_0_control_slave_readdata
	wire    [2:0] mm_interconnect_2_performance_counter_0_control_slave_address;                // mm_interconnect_2:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire          mm_interconnect_2_performance_counter_0_control_slave_begintransfer;          // mm_interconnect_2:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire          mm_interconnect_2_performance_counter_0_control_slave_write;                  // mm_interconnect_2:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire   [31:0] mm_interconnect_2_performance_counter_0_control_slave_writedata;              // mm_interconnect_2:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire   [31:0] mm_interconnect_2_msgdma_0_csr_readdata;                                      // msgdma_0:csr_readdata -> mm_interconnect_2:msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_2_msgdma_0_csr_address;                                       // mm_interconnect_2:msgdma_0_csr_address -> msgdma_0:csr_address
	wire          mm_interconnect_2_msgdma_0_csr_read;                                          // mm_interconnect_2:msgdma_0_csr_read -> msgdma_0:csr_read
	wire    [3:0] mm_interconnect_2_msgdma_0_csr_byteenable;                                    // mm_interconnect_2:msgdma_0_csr_byteenable -> msgdma_0:csr_byteenable
	wire          mm_interconnect_2_msgdma_0_csr_write;                                         // mm_interconnect_2:msgdma_0_csr_write -> msgdma_0:csr_write
	wire   [31:0] mm_interconnect_2_msgdma_0_csr_writedata;                                     // mm_interconnect_2:msgdma_0_csr_writedata -> msgdma_0:csr_writedata
	wire   [31:0] mm_interconnect_2_vic_0_csr_access_readdata;                                  // vic_0:csr_access_readdata -> mm_interconnect_2:vic_0_csr_access_readdata
	wire    [7:0] mm_interconnect_2_vic_0_csr_access_address;                                   // mm_interconnect_2:vic_0_csr_access_address -> vic_0:csr_access_address
	wire          mm_interconnect_2_vic_0_csr_access_read;                                      // mm_interconnect_2:vic_0_csr_access_read -> vic_0:csr_access_read
	wire          mm_interconnect_2_vic_0_csr_access_write;                                     // mm_interconnect_2:vic_0_csr_access_write -> vic_0:csr_access_write
	wire   [31:0] mm_interconnect_2_vic_0_csr_access_writedata;                                 // mm_interconnect_2:vic_0_csr_access_writedata -> vic_0:csr_access_writedata
	wire          mm_interconnect_2_msgdma_0_descriptor_slave_waitrequest;                      // msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_2:msgdma_0_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_2_msgdma_0_descriptor_slave_byteenable;                       // mm_interconnect_2:msgdma_0_descriptor_slave_byteenable -> msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_2_msgdma_0_descriptor_slave_write;                            // mm_interconnect_2:msgdma_0_descriptor_slave_write -> msgdma_0:descriptor_slave_write
	wire  [127:0] mm_interconnect_2_msgdma_0_descriptor_slave_writedata;                        // mm_interconnect_2:msgdma_0_descriptor_slave_writedata -> msgdma_0:descriptor_slave_writedata
	wire          mm_interconnect_2_timer_0_s1_chipselect;                                      // mm_interconnect_2:timer_0_s1_chipselect -> timer_0:chipselect
	wire   [15:0] mm_interconnect_2_timer_0_s1_readdata;                                        // timer_0:readdata -> mm_interconnect_2:timer_0_s1_readdata
	wire    [2:0] mm_interconnect_2_timer_0_s1_address;                                         // mm_interconnect_2:timer_0_s1_address -> timer_0:address
	wire          mm_interconnect_2_timer_0_s1_write;                                           // mm_interconnect_2:timer_0_s1_write -> timer_0:write_n
	wire   [15:0] mm_interconnect_2_timer_0_s1_writedata;                                       // mm_interconnect_2:timer_0_s1_writedata -> timer_0:writedata
	wire          mm_bridge_1_m0_waitrequest;                                                   // mm_interconnect_3:mm_bridge_1_m0_waitrequest -> mm_bridge_1:m0_waitrequest
	wire   [31:0] mm_bridge_1_m0_readdata;                                                      // mm_interconnect_3:mm_bridge_1_m0_readdata -> mm_bridge_1:m0_readdata
	wire          mm_bridge_1_m0_debugaccess;                                                   // mm_bridge_1:m0_debugaccess -> mm_interconnect_3:mm_bridge_1_m0_debugaccess
	wire   [12:0] mm_bridge_1_m0_address;                                                       // mm_bridge_1:m0_address -> mm_interconnect_3:mm_bridge_1_m0_address
	wire          mm_bridge_1_m0_read;                                                          // mm_bridge_1:m0_read -> mm_interconnect_3:mm_bridge_1_m0_read
	wire    [3:0] mm_bridge_1_m0_byteenable;                                                    // mm_bridge_1:m0_byteenable -> mm_interconnect_3:mm_bridge_1_m0_byteenable
	wire          mm_bridge_1_m0_readdatavalid;                                                 // mm_interconnect_3:mm_bridge_1_m0_readdatavalid -> mm_bridge_1:m0_readdatavalid
	wire   [31:0] mm_bridge_1_m0_writedata;                                                     // mm_bridge_1:m0_writedata -> mm_interconnect_3:mm_bridge_1_m0_writedata
	wire          mm_bridge_1_m0_write;                                                         // mm_bridge_1:m0_write -> mm_interconnect_3:mm_bridge_1_m0_write
	wire    [0:0] mm_bridge_1_m0_burstcount;                                                    // mm_bridge_1:m0_burstcount -> mm_interconnect_3:mm_bridge_1_m0_burstcount
	wire          mm_interconnect_3_pio_0_s1_chipselect;                                        // mm_interconnect_3:pio_0_s1_chipselect -> pio_0:chipselect
	wire   [31:0] mm_interconnect_3_pio_0_s1_readdata;                                          // pio_0:readdata -> mm_interconnect_3:pio_0_s1_readdata
	wire    [1:0] mm_interconnect_3_pio_0_s1_address;                                           // mm_interconnect_3:pio_0_s1_address -> pio_0:address
	wire          mm_interconnect_3_pio_0_s1_write;                                             // mm_interconnect_3:pio_0_s1_write -> pio_0:write_n
	wire   [31:0] mm_interconnect_3_pio_0_s1_writedata;                                         // mm_interconnect_3:pio_0_s1_writedata -> pio_0:writedata
	wire          mm_interconnect_3_pio_1_s1_chipselect;                                        // mm_interconnect_3:pio_1_s1_chipselect -> pio_1:chipselect
	wire   [31:0] mm_interconnect_3_pio_1_s1_readdata;                                          // pio_1:readdata -> mm_interconnect_3:pio_1_s1_readdata
	wire    [1:0] mm_interconnect_3_pio_1_s1_address;                                           // mm_interconnect_3:pio_1_s1_address -> pio_1:address
	wire          mm_interconnect_3_pio_1_s1_write;                                             // mm_interconnect_3:pio_1_s1_write -> pio_1:write_n
	wire   [31:0] mm_interconnect_3_pio_1_s1_writedata;                                         // mm_interconnect_3:pio_1_s1_writedata -> pio_1:writedata
	wire          mm_interconnect_3_pio_2_s1_chipselect;                                        // mm_interconnect_3:pio_2_s1_chipselect -> pio_2:chipselect
	wire   [31:0] mm_interconnect_3_pio_2_s1_readdata;                                          // pio_2:readdata -> mm_interconnect_3:pio_2_s1_readdata
	wire    [2:0] mm_interconnect_3_pio_2_s1_address;                                           // mm_interconnect_3:pio_2_s1_address -> pio_2:address
	wire          mm_interconnect_3_pio_2_s1_write;                                             // mm_interconnect_3:pio_2_s1_write -> pio_2:write_n
	wire   [31:0] mm_interconnect_3_pio_2_s1_writedata;                                         // mm_interconnect_3:pio_2_s1_writedata -> pio_2:writedata
	wire   [15:0] mm_interconnect_3_motor_controller_5_slave_readdata;                          // motor_controller_5:slave_readdata -> mm_interconnect_3:motor_controller_5_slave_readdata
	wire    [1:0] mm_interconnect_3_motor_controller_5_slave_address;                           // mm_interconnect_3:motor_controller_5_slave_address -> motor_controller_5:slave_address
	wire          mm_interconnect_3_motor_controller_5_slave_read;                              // mm_interconnect_3:motor_controller_5_slave_read -> motor_controller_5:slave_read
	wire          mm_interconnect_3_motor_controller_5_slave_write;                             // mm_interconnect_3:motor_controller_5_slave_write -> motor_controller_5:slave_write
	wire   [15:0] mm_interconnect_3_motor_controller_5_slave_writedata;                         // mm_interconnect_3:motor_controller_5_slave_writedata -> motor_controller_5:slave_writedata
	wire   [15:0] mm_interconnect_3_imu_spim_slave_readdata;                                    // imu_spim:slave_readdata -> mm_interconnect_3:imu_spim_slave_readdata
	wire    [2:0] mm_interconnect_3_imu_spim_slave_address;                                     // mm_interconnect_3:imu_spim_slave_address -> imu_spim:slave_address
	wire          mm_interconnect_3_imu_spim_slave_read;                                        // mm_interconnect_3:imu_spim_slave_read -> imu_spim:slave_read
	wire          mm_interconnect_3_imu_spim_slave_write;                                       // mm_interconnect_3:imu_spim_slave_write -> imu_spim:slave_write
	wire   [15:0] mm_interconnect_3_imu_spim_slave_writedata;                                   // mm_interconnect_3:imu_spim_slave_writedata -> imu_spim:slave_writedata
	wire   [15:0] mm_interconnect_3_i2c_master_0_slave_readdata;                                // i2c_master_0:slave_readdata -> mm_interconnect_3:i2c_master_0_slave_readdata
	wire    [2:0] mm_interconnect_3_i2c_master_0_slave_address;                                 // mm_interconnect_3:i2c_master_0_slave_address -> i2c_master_0:slave_address
	wire          mm_interconnect_3_i2c_master_0_slave_read;                                    // mm_interconnect_3:i2c_master_0_slave_read -> i2c_master_0:slave_read
	wire          mm_interconnect_3_i2c_master_0_slave_write;                                   // mm_interconnect_3:i2c_master_0_slave_write -> i2c_master_0:slave_write
	wire   [15:0] mm_interconnect_3_i2c_master_0_slave_writedata;                               // mm_interconnect_3:i2c_master_0_slave_writedata -> i2c_master_0:slave_writedata
	wire   [15:0] mm_interconnect_3_vector_controller_master_0_slave_readdata;                  // vector_controller_master_0:slave_readdata -> mm_interconnect_3:vector_controller_master_0_slave_readdata
	wire    [4:0] mm_interconnect_3_vector_controller_master_0_slave_address;                   // mm_interconnect_3:vector_controller_master_0_slave_address -> vector_controller_master_0:slave_address
	wire          mm_interconnect_3_vector_controller_master_0_slave_read;                      // mm_interconnect_3:vector_controller_master_0_slave_read -> vector_controller_master_0:slave_read
	wire          mm_interconnect_3_vector_controller_master_0_slave_write;                     // mm_interconnect_3:vector_controller_master_0_slave_write -> vector_controller_master_0:slave_write
	wire   [15:0] mm_interconnect_3_vector_controller_master_0_slave_writedata;                 // mm_interconnect_3:vector_controller_master_0_slave_writedata -> vector_controller_master_0:slave_writedata
	wire          mm_interconnect_3_spim_0_spi_control_port_chipselect;                         // mm_interconnect_3:spim_0_spi_control_port_chipselect -> spim_0:spi_select
	wire   [15:0] mm_interconnect_3_spim_0_spi_control_port_readdata;                           // spim_0:data_to_cpu -> mm_interconnect_3:spim_0_spi_control_port_readdata
	wire    [2:0] mm_interconnect_3_spim_0_spi_control_port_address;                            // mm_interconnect_3:spim_0_spi_control_port_address -> spim_0:mem_addr
	wire          mm_interconnect_3_spim_0_spi_control_port_read;                               // mm_interconnect_3:spim_0_spi_control_port_read -> spim_0:read_n
	wire          mm_interconnect_3_spim_0_spi_control_port_write;                              // mm_interconnect_3:spim_0_spi_control_port_write -> spim_0:write_n
	wire   [15:0] mm_interconnect_3_spim_0_spi_control_port_writedata;                          // mm_interconnect_3:spim_0_spi_control_port_writedata -> spim_0:data_from_cpu
	wire          mm_bridge_2_m0_waitrequest;                                                   // mm_interconnect_4:mm_bridge_2_m0_waitrequest -> mm_bridge_2:m0_waitrequest
	wire   [31:0] mm_bridge_2_m0_readdata;                                                      // mm_interconnect_4:mm_bridge_2_m0_readdata -> mm_bridge_2:m0_readdata
	wire          mm_bridge_2_m0_debugaccess;                                                   // mm_bridge_2:m0_debugaccess -> mm_interconnect_4:mm_bridge_2_m0_debugaccess
	wire   [14:0] mm_bridge_2_m0_address;                                                       // mm_bridge_2:m0_address -> mm_interconnect_4:mm_bridge_2_m0_address
	wire          mm_bridge_2_m0_read;                                                          // mm_bridge_2:m0_read -> mm_interconnect_4:mm_bridge_2_m0_read
	wire    [3:0] mm_bridge_2_m0_byteenable;                                                    // mm_bridge_2:m0_byteenable -> mm_interconnect_4:mm_bridge_2_m0_byteenable
	wire          mm_bridge_2_m0_readdatavalid;                                                 // mm_interconnect_4:mm_bridge_2_m0_readdatavalid -> mm_bridge_2:m0_readdatavalid
	wire   [31:0] mm_bridge_2_m0_writedata;                                                     // mm_bridge_2:m0_writedata -> mm_interconnect_4:mm_bridge_2_m0_writedata
	wire          mm_bridge_2_m0_write;                                                         // mm_bridge_2:m0_write -> mm_interconnect_4:mm_bridge_2_m0_write
	wire    [0:0] mm_bridge_2_m0_burstcount;                                                    // mm_bridge_2:m0_burstcount -> mm_interconnect_4:mm_bridge_2_m0_burstcount
	wire    [7:0] msgdma_0_mm_read_readdata;                                                    // mm_interconnect_4:msgdma_0_mm_read_readdata -> msgdma_0:mm_read_readdata
	wire          msgdma_0_mm_read_waitrequest;                                                 // mm_interconnect_4:msgdma_0_mm_read_waitrequest -> msgdma_0:mm_read_waitrequest
	wire   [15:0] msgdma_0_mm_read_address;                                                     // msgdma_0:mm_read_address -> mm_interconnect_4:msgdma_0_mm_read_address
	wire          msgdma_0_mm_read_read;                                                        // msgdma_0:mm_read_read -> mm_interconnect_4:msgdma_0_mm_read_read
	wire          msgdma_0_mm_read_readdatavalid;                                               // mm_interconnect_4:msgdma_0_mm_read_readdatavalid -> msgdma_0:mm_read_readdatavalid
	wire          mm_interconnect_4_instruction_rom_0_s2_chipselect;                            // mm_interconnect_4:instruction_rom_0_s2_chipselect -> instruction_rom_0:chipselect2
	wire   [31:0] mm_interconnect_4_instruction_rom_0_s2_readdata;                              // instruction_rom_0:readdata2 -> mm_interconnect_4:instruction_rom_0_s2_readdata
	wire   [12:0] mm_interconnect_4_instruction_rom_0_s2_address;                               // mm_interconnect_4:instruction_rom_0_s2_address -> instruction_rom_0:address2
	wire    [3:0] mm_interconnect_4_instruction_rom_0_s2_byteenable;                            // mm_interconnect_4:instruction_rom_0_s2_byteenable -> instruction_rom_0:byteenable2
	wire          mm_interconnect_4_instruction_rom_0_s2_write;                                 // mm_interconnect_4:instruction_rom_0_s2_write -> instruction_rom_0:write2
	wire   [31:0] mm_interconnect_4_instruction_rom_0_s2_writedata;                             // mm_interconnect_4:instruction_rom_0_s2_writedata -> instruction_rom_0:writedata2
	wire          mm_interconnect_4_instruction_rom_0_s2_clken;                                 // mm_interconnect_4:instruction_rom_0_s2_clken -> instruction_rom_0:clken2
	wire          mm_interconnect_4_data_ram_0_s2_chipselect;                                   // mm_interconnect_4:data_ram_0_s2_chipselect -> data_ram_0:chipselect2
	wire   [31:0] mm_interconnect_4_data_ram_0_s2_readdata;                                     // data_ram_0:readdata2 -> mm_interconnect_4:data_ram_0_s2_readdata
	wire    [9:0] mm_interconnect_4_data_ram_0_s2_address;                                      // mm_interconnect_4:data_ram_0_s2_address -> data_ram_0:address2
	wire    [3:0] mm_interconnect_4_data_ram_0_s2_byteenable;                                   // mm_interconnect_4:data_ram_0_s2_byteenable -> data_ram_0:byteenable2
	wire          mm_interconnect_4_data_ram_0_s2_write;                                        // mm_interconnect_4:data_ram_0_s2_write -> data_ram_0:write2
	wire   [31:0] mm_interconnect_4_data_ram_0_s2_writedata;                                    // mm_interconnect_4:data_ram_0_s2_writedata -> data_ram_0:writedata2
	wire          mm_interconnect_4_data_ram_0_s2_clken;                                        // mm_interconnect_4:data_ram_0_s2_clken -> data_ram_0:clken2
	wire          irq_mapper_receiver0_irq;                                                     // msgdma_0:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                     // spim_0:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                     // pio_0:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                     // pio_1:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                     // vector_controller_master_0:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                     // motor_controller_5:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                     // timer_0:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                     // i2c_master_0:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                     // jtag_uart_0:av_irq -> irq_mapper:receiver8_irq
	wire    [8:0] vic_0_irq_input_irq;                                                          // irq_mapper:sender_irq -> vic_0:irq_input_irq
	wire          rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [data_ram_0:reset, data_ram_1:reset, instruction_rom_0:reset, mm_bridge_2:reset, mm_interconnect_0:spi_slave_to_avalon_mm_master_bridge_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:instruction_rom_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_4:mm_bridge_2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, spi_slave_to_avalon_mm_master_bridge_0:reset_n]
	wire          rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [data_ram_0:reset_req, data_ram_1:reset_req, instruction_rom_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                           // rst_controller_001:reset_out -> [dc_fifo_0:in_reset_n, i2c_master_0:reset, imu_spim:reset, irq_mapper:reset, mm_bridge_1:reset, mm_interconnect_1:mm_bridge_1_reset_reset_bridge_in_reset_reset, mm_interconnect_2:performance_counter_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:mm_bridge_1_reset_reset_bridge_in_reset_reset, mm_interconnect_3:motor_controller_5_reset_reset_bridge_in_reset_reset, mm_interconnect_4:msgdma_0_reset_n_reset_bridge_in_reset_reset, msgdma_0:reset_n_reset_n, performance_counter_0:reset_n, pio_0:reset_n, pio_1:reset_n, pio_2:reset_n, spim_0:reset_n, st_packets_to_bytes_0:reset_n, timer_0:reset_n, vector_controller_master_0:reset, vic_0:reset_reset]
	wire          nios_0_debug_reset_request_reset;                                             // nios_0:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_004:reset_in1]
	wire          reset_controller_0_reset_out_reset;                                           // reset_controller_0:reset_out -> [rst_controller_001:reset_in2, rst_controller_003:reset_in1, rst_controller_004:reset_in2]
	wire          rst_controller_002_reset_out_reset;                                           // rst_controller_002:reset_out -> dc_fifo_0:out_reset_n
	wire          rst_controller_003_reset_out_reset;                                           // rst_controller_003:reset_out -> [jtag_uart_0:rst_n, mm_bridge_0:reset, mm_interconnect_1:nios_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_bridge_0_reset_reset_bridge_in_reset_reset, nios_0:reset_n, rst_translator_001:in_reset, sysid_qsys_0:reset_n]
	wire          rst_controller_003_reset_out_reset_req;                                       // rst_controller_003:reset_req -> [nios_0:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_004_reset_out_reset;                                           // rst_controller_004:reset_out -> motor_controller_5:reset

	avalon_st_uart_tx #(
		.PRESCALER (25)
	) avalon_st_uart_tx_0 (
		.clk        (clk_100mhz_clk),        //   clk.clk
		.reset      (~reset_100mhz_reset_n), // reset.reset
		.sink_ready (dc_fifo_0_out_ready),   //  sink.ready
		.sink_valid (dc_fifo_0_out_valid),   //      .valid
		.sink_data  (dc_fifo_0_out_data),    //      .data
		.uart_txd   (uart_txd)               //  uart.txd
	);

	controller_data_ram_0 data_ram_0 (
		.address     (mm_interconnect_1_data_ram_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_data_ram_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_data_ram_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_data_ram_0_s1_write),      //       .write
		.readdata    (mm_interconnect_1_data_ram_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_data_ram_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_data_ram_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_4_data_ram_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_4_data_ram_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_4_data_ram_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_4_data_ram_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_4_data_ram_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_4_data_ram_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_4_data_ram_0_s2_byteenable), //       .byteenable
		.clk         (clk_sys_clk),                                //   clk1.clk
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	controller_data_ram_1 data_ram_1 (
		.address     (mm_interconnect_1_data_ram_1_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_data_ram_1_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_data_ram_1_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_data_ram_1_s1_write),      //       .write
		.readdata    (mm_interconnect_1_data_ram_1_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_data_ram_1_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_data_ram_1_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_data_ram_1_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_data_ram_1_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_data_ram_1_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_data_ram_1_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_data_ram_1_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_data_ram_1_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_data_ram_1_s2_byteenable), //       .byteenable
		.clk         (clk_sys_clk),                                //   clk1.clk
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (8),
		.FIFO_DEPTH         (128),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dc_fifo_0 (
		.in_clk            (clk_sys_clk),                                  //        in_clk.clk
		.in_reset_n        (~rst_controller_001_reset_out_reset),          //  in_clk_reset.reset_n
		.out_clk           (clk_100mhz_clk),                               //       out_clk.clk
		.out_reset_n       (~rst_controller_002_reset_out_reset),          // out_clk_reset.reset_n
		.in_data           (st_packets_to_bytes_0_out_bytes_stream_data),  //            in.data
		.in_valid          (st_packets_to_bytes_0_out_bytes_stream_valid), //              .valid
		.in_ready          (st_packets_to_bytes_0_out_bytes_stream_ready), //              .ready
		.out_data          (dc_fifo_0_out_data),                           //           out.data
		.out_valid         (dc_fifo_0_out_valid),                          //              .valid
		.out_ready         (dc_fifo_0_out_ready),                          //              .ready
		.in_csr_address    (1'b0),                                         //   (terminated)
		.in_csr_read       (1'b0),                                         //   (terminated)
		.in_csr_write      (1'b0),                                         //   (terminated)
		.in_csr_readdata   (),                                             //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000),         //   (terminated)
		.out_csr_address   (1'b0),                                         //   (terminated)
		.out_csr_read      (1'b0),                                         //   (terminated)
		.out_csr_write     (1'b0),                                         //   (terminated)
		.out_csr_readdata  (),                                             //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000),         //   (terminated)
		.in_startofpacket  (1'b0),                                         //   (terminated)
		.in_endofpacket    (1'b0),                                         //   (terminated)
		.out_startofpacket (),                                             //   (terminated)
		.out_endofpacket   (),                                             //   (terminated)
		.in_empty          (1'b0),                                         //   (terminated)
		.out_empty         (),                                             //   (terminated)
		.in_error          (1'b0),                                         //   (terminated)
		.out_error         (),                                             //   (terminated)
		.in_channel        (1'b0),                                         //   (terminated)
		.out_channel       (),                                             //   (terminated)
		.space_avail_data  ()                                              //   (terminated)
	);

	float32to16 float32to16_0 (
		.slave_reset  (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  // slave.reset
		.slave_clk    (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //      .clk
		.slave_clk_en (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //      .clk_en
		.slave_start  (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //      .start
		.slave_done   (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //      .done
		.slave_dataa  (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //      .dataa
		.slave_result (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_result)  //      .result
	);

	controller_fpu_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) fpu_0 (
		.s1_dataa     (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),       // s2.clk
		.s2_clk_en    (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),     //   .dataa
		.s2_datab     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),     //   .datab
		.s2_n         (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_n),         //   .n
		.s2_reset     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),     //   .reset
		.s2_reset_req (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset_req), //   .reset_req
		.s2_start     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_start),     //   .start
		.s2_done      (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_done),      //   .done
		.s2_result    (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_result)     //   .result
	);

	i2c_master #(
		.PRESCALER (188)
	) i2c_master_0 (
		.clk             (clk_sys_clk),                                    //   clk.clk
		.reset           (rst_controller_001_reset_out_reset),             // reset.reset
		.slave_address   (mm_interconnect_3_i2c_master_0_slave_address),   // slave.address
		.slave_read      (mm_interconnect_3_i2c_master_0_slave_read),      //      .read
		.slave_readdata  (mm_interconnect_3_i2c_master_0_slave_readdata),  //      .readdata
		.slave_write     (mm_interconnect_3_i2c_master_0_slave_write),     //      .write
		.slave_writedata (mm_interconnect_3_i2c_master_0_slave_writedata), //      .writedata
		.irq             (irq_mapper_receiver7_irq),                       //   irq.irq
		.i2c_scl_in      (adc2_i2c_scl_in),                                //   i2c.scl_in
		.i2c_sda_in      (adc2_i2c_sda_in),                                //      .sda_in
		.i2c_scl_oe      (adc2_i2c_scl_oe),                                //      .scl_oe
		.i2c_sda_oe      (adc2_i2c_sda_oe)                                 //      .sda_oe
	);

	imu_spim #(
		.PRESCALER (2)
	) imu_spim (
		.reset           (rst_controller_001_reset_out_reset),         // reset.reset
		.clk             (clk_sys_clk),                                //   clk.clk
		.slave_address   (mm_interconnect_3_imu_spim_slave_address),   // slave.address
		.slave_read      (mm_interconnect_3_imu_spim_slave_read),      //      .read
		.slave_readdata  (mm_interconnect_3_imu_spim_slave_readdata),  //      .readdata
		.slave_write     (mm_interconnect_3_imu_spim_slave_write),     //      .write
		.slave_writedata (mm_interconnect_3_imu_spim_slave_writedata), //      .writedata
		.SCLK            (spim_0_external_sclk),                       //  spis.export
		.MOSI            (spim_0_external_mosi),                       //      .export
		.MISO            (imu_spim_spis_miso),                         //      .export
		.SS_n            (spim_0_external_ss_n),                       //      .export
		.spim_mosi       (imu_spi_mosi),                               //  spim.mosi
		.spim_miso       (imu_spi_miso),                               //      .miso
		.spim_sclk       (imu_spi_sclk),                               //      .sclk
		.spim_cs_n       (imu_spi_cs_n),                               //      .cs_n
		.spim_int_n      (imu_spi_int_n)                               //      .int_n
	);

	controller_instruction_rom_0 instruction_rom_0 (
		.address     (mm_interconnect_1_instruction_rom_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_instruction_rom_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_instruction_rom_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_instruction_rom_0_s1_write),      //       .write
		.readdata    (mm_interconnect_1_instruction_rom_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_instruction_rom_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_instruction_rom_0_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_4_instruction_rom_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_4_instruction_rom_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_4_instruction_rom_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_4_instruction_rom_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_4_instruction_rom_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_4_instruction_rom_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_4_instruction_rom_0_s2_byteenable), //       .byteenable
		.clk         (clk_sys_clk),                                       //   clk1.clk
		.reset       (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze      (1'b0)                                               // (terminated)
	);

	controller_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_sys_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver8_irq)                                     //               irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_sys_clk),                                    //   clk.clk
		.reset            (rst_controller_003_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (13),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_1 (
		.clk              (clk_sys_clk),                                    //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_1_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_1_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_1_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_1_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_1_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_1_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_1_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_1_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_1_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_1_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_1_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_1_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_1_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_1_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_1_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_1_m0_address),                         //      .address
		.m0_write         (mm_bridge_1_m0_write),                           //      .write
		.m0_read          (mm_bridge_1_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_1_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_1_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (15),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_2 (
		.clk              (clk_sys_clk),                                    //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_2_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_2_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_2_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_2_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_2_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_2_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_2_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_2_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_2_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_2_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_2_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_2_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_2_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_2_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_2_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_2_m0_address),                         //      .address
		.m0_write         (mm_bridge_2_m0_write),                           //      .write
		.m0_read          (mm_bridge_2_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_2_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_2_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                               // (terminated)
		.m0_response      (2'b00)                                           // (terminated)
	);

	motor_controller motor_controller_5 (
		.clk                   (clk_sys_clk),                                          //        clk.clk
		.reset                 (rst_controller_004_reset_out_reset),                   //      reset.reset
		.fault                 (mc5_fault_fault),                                      //      fault.fault
		.brake                 (mc5_fault_brake),                                      //           .brake
		.status_driver_otw_n   (mc5_status_driver_otw_n),                              //     status.driver_otw_n
		.status_driver_fault_n (mc5_status_driver_fault_n),                            //           .driver_fault_n
		.status_hall_fault_n   (mc5_status_hall_fault_n),                              //           .hall_fault_n
		.pwm_source_data       (mc5_pwm_data),                                         // pwm_source.data
		.pwm_source_valid      (mc5_pwm_valid),                                        //           .valid
		.pwm_source_ready      (mc5_pwm_ready),                                        //           .ready
		.slave_address         (mm_interconnect_3_motor_controller_5_slave_address),   //      slave.address
		.slave_readdata        (mm_interconnect_3_motor_controller_5_slave_readdata),  //           .readdata
		.slave_writedata       (mm_interconnect_3_motor_controller_5_slave_writedata), //           .writedata
		.slave_read            (mm_interconnect_3_motor_controller_5_slave_read),      //           .read
		.slave_write           (mm_interconnect_3_motor_controller_5_slave_write),     //           .write
		.irq                   (irq_mapper_receiver5_irq)                              //        irq.irq
	);

	controller_msgdma_0 msgdma_0 (
		.mm_read_address              (msgdma_0_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (msgdma_0_mm_read_read),                                   //                 .read
		.mm_read_readdata             (msgdma_0_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (msgdma_0_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (msgdma_0_mm_read_readdatavalid),                          //                 .readdatavalid
		.clock_clk                    (clk_sys_clk),                                             //            clock.clk
		.reset_n_reset_n              (~rst_controller_001_reset_out_reset),                     //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_2_msgdma_0_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_2_msgdma_0_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_2_msgdma_0_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_2_msgdma_0_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_2_msgdma_0_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_2_msgdma_0_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_2_msgdma_0_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_2_msgdma_0_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_2_msgdma_0_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_2_msgdma_0_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                //          csr_irq.irq
		.st_source_data               (msgdma_0_st_source_data),                                 //        st_source.data
		.st_source_valid              (msgdma_0_st_source_valid),                                //                 .valid
		.st_source_ready              (msgdma_0_st_source_ready),                                //                 .ready
		.st_source_startofpacket      (msgdma_0_st_source_startofpacket),                        //                 .startofpacket
		.st_source_endofpacket        (msgdma_0_st_source_endofpacket),                          //                 .endofpacket
		.st_source_channel            (msgdma_0_st_source_channel)                               //                 .channel
	);

	controller_nios_0 nios_0 (
		.clk                                 (clk_sys_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),               //                          .reset_req
		.d_address                           (nios_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_0_data_master_read),                              //                          .read
		.d_readdata                          (nios_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_0_data_master_write),                             //                          .write
		.d_writedata                         (nios_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_0_instruction_master_waitrequest),                //                          .waitrequest
		.eic_port_valid                      (vic_0_interrupt_controller_out_valid),                 //   interrupt_controller_in.valid
		.eic_port_data                       (vic_0_interrupt_controller_out_data),                  //                          .data
		.debug_reset_request                 (nios_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios_0_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios_0_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios_0_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios_0_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios_0_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios_0_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios_0_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios_0_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios_0_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios_0_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios_0_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios_0_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios_0_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios_0_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios_0_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios_0_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios_0_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (nios_0_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (nios_0_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (nios_0_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (nios_0_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (nios_0_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (nios_0_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (nios_0_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (nios_0_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (nios_0_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (nios_0_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (nios_0_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (nios_0_custom_instruction_master_writerc)              //                          .writerc
	);

	controller_performance_counter_0 performance_counter_0 (
		.clk           (clk_sys_clk),                                                         //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                                 //         reset.reset_n
		.address       (mm_interconnect_2_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_2_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_2_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_2_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_2_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	controller_pio_0 pio_0 (
		.clk        (clk_sys_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_3_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_pio_0_s1_readdata),   //                    .readdata
		.in_port    (pio_0_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)               //                 irq.irq
	);

	controller_pio_1 pio_1 (
		.clk        (clk_sys_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_3_pio_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_pio_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_pio_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_pio_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_pio_1_s1_readdata),   //                    .readdata
		.in_port    (pio_1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)               //                 irq.irq
	);

	controller_pio_2 pio_2 (
		.clk        (clk_sys_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_3_pio_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_pio_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_pio_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_pio_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_pio_2_s1_readdata),   //                    .readdata
		.out_port   (pio_2_export)                           // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_0 (
		.reset_in0      (reset_ext_reset),                    // reset_in0.reset
		.clk            (clk_sys_clk),                        //       clk.clk
		.reset_out      (reset_controller_0_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	SPISlaveToAvalonMasterBridge #(
		.SYNC_DEPTH (2)
	) spi_slave_to_avalon_mm_master_bridge_0 (
		.clk                                                                    (clk_sys_clk),                                                        //           clk.clk
		.reset_n                                                                (~rst_controller_reset_out_reset),                                    //     clk_reset.reset_n
		.mosi_to_the_spislave_inst_for_spichain                                 (host_spi_mosi_to_the_spislave_inst_for_spichain),                    //      export_0.export
		.nss_to_the_spislave_inst_for_spichain                                  (host_spi_nss_to_the_spislave_inst_for_spichain),                     //              .export
		.miso_to_and_from_the_spislave_inst_for_spichain                        (host_spi_miso_to_and_from_the_spislave_inst_for_spichain),           //              .export
		.sclk_to_the_spislave_inst_for_spichain                                 (host_spi_sclk_to_the_spislave_inst_for_spichain),                    //              .export
		.address_from_the_altera_avalon_packets_to_master_inst_for_spichain     (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address),       // avalon_master.address
		.byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain  (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable),    //              .byteenable
		.read_from_the_altera_avalon_packets_to_master_inst_for_spichain        (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read),          //              .read
		.readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain      (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata),      //              .readdata
		.readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid), //              .readdatavalid
		.waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest),   //              .waitrequest
		.write_from_the_altera_avalon_packets_to_master_inst_for_spichain       (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write),         //              .write
		.writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata)      //              .writedata
	);

	controller_spim_0 spim_0 (
		.clk           (clk_sys_clk),                                          //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                  //            reset.reset_n
		.data_from_cpu (mm_interconnect_3_spim_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_3_spim_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_3_spim_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_3_spim_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_3_spim_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_3_spim_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                             //              irq.irq
		.MISO          (imu_spim_spis_miso),                                   //         external.export
		.MOSI          (spim_0_external_mosi),                                 //                 .export
		.SCLK          (spim_0_external_sclk),                                 //                 .export
		.SS_n          (spim_0_external_ss_n)                                  //                 .export
	);

	altera_avalon_st_packets_to_bytes #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_packets_to_bytes_0 (
		.clk              (clk_sys_clk),                                  //               clk.clk
		.reset_n          (~rst_controller_001_reset_out_reset),          //         clk_reset.reset_n
		.in_ready         (msgdma_0_st_source_ready),                     // in_packets_stream.ready
		.in_valid         (msgdma_0_st_source_valid),                     //                  .valid
		.in_data          (msgdma_0_st_source_data),                      //                  .data
		.in_channel       (msgdma_0_st_source_channel),                   //                  .channel
		.in_startofpacket (msgdma_0_st_source_startofpacket),             //                  .startofpacket
		.in_endofpacket   (msgdma_0_st_source_endofpacket),               //                  .endofpacket
		.out_ready        (st_packets_to_bytes_0_out_bytes_stream_ready), //  out_bytes_stream.ready
		.out_valid        (st_packets_to_bytes_0_out_bytes_stream_valid), //                  .valid
		.out_data         (st_packets_to_bytes_0_out_bytes_stream_data)   //                  .data
	);

	controller_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_sys_clk),                                           //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_0_control_slave_address)   //              .address
	);

	controller_timer_0 timer_0 (
		.clk        (clk_sys_clk),                             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_2_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_2_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_2_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_2_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_2_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver6_irq)                 //   irq.irq
	);

	vector_controller_master vector_controller_master_0 (
		.clk                         (clk_sys_clk),                                                  //                   clk.clk
		.reset                       (rst_controller_001_reset_out_reset),                           //                 reset.reset
		.fault                       (vc_fault_fault),                                               //                 fault.fault
		.brake                       (vc_fault_brake),                                               //                      .brake
		.status_driver_otw_n         (vc_status_driver_otw_n),                                       //                status.driver_otw_n
		.status_driver_fault_n       (vc_status_driver_fault_n),                                     //                      .driver_fault_n
		.status_hall_fault_n         (vc_status_hall_fault_n),                                       //                      .hall_fault_n
		.status_encoder_fault_n      (vc_status_encoder_fault_n),                                    //                      .encoder_fault_n
		.status_pos_error            (vc_status_pos_error),                                          //                      .pos_error
		.status_pos_uncertain        (vc_status_pos_uncertain),                                      //                      .pos_uncertain
		.encoder_1_data              (vc_encoder_encoder_1_data),                                    //               encoder.encoder_1_data
		.encoder_2_data              (vc_encoder_encoder_2_data),                                    //                      .encoder_2_data
		.encoder_3_data              (vc_encoder_encoder_3_data),                                    //                      .encoder_3_data
		.encoder_4_data              (vc_encoder_encoder_4_data),                                    //                      .encoder_4_data
		.param_kp                    (vc_param_kp),                                                  //                 param.kp
		.param_ki                    (vc_param_ki),                                                  //                      .ki
		.current_measurement_1_data  (vc_imeas1_data),                                               // current_measurement_1.data
		.current_measurement_1_valid (vc_imeas1_valid),                                              //                      .valid
		.current_measurement_2_data  (vc_imeas2_data),                                               // current_measurement_2.data
		.current_measurement_2_valid (vc_imeas2_valid),                                              //                      .valid
		.current_measurement_3_data  (vc_imeas3_data),                                               // current_measurement_3.data
		.current_measurement_3_valid (vc_imeas3_valid),                                              //                      .valid
		.current_measurement_4_data  (vc_imeas4_data),                                               // current_measurement_4.data
		.current_measurement_4_valid (vc_imeas4_valid),                                              //                      .valid
		.current_reference_1_data    (vc_iref1_data),                                                //   current_reference_1.data
		.current_reference_1_valid   (vc_iref1_valid),                                               //                      .valid
		.current_reference_2_data    (vc_iref2_data),                                                //   current_reference_2.data
		.current_reference_2_valid   (vc_iref2_valid),                                               //                      .valid
		.current_reference_3_data    (vc_iref3_data),                                                //   current_reference_3.data
		.current_reference_3_valid   (vc_iref3_valid),                                               //                      .valid
		.current_reference_4_data    (vc_iref4_data),                                                //   current_reference_4.data
		.current_reference_4_valid   (vc_iref4_valid),                                               //                      .valid
		.slave_address               (mm_interconnect_3_vector_controller_master_0_slave_address),   //                 slave.address
		.slave_read                  (mm_interconnect_3_vector_controller_master_0_slave_read),      //                      .read
		.slave_readdata              (mm_interconnect_3_vector_controller_master_0_slave_readdata),  //                      .readdata
		.slave_write                 (mm_interconnect_3_vector_controller_master_0_slave_write),     //                      .write
		.slave_writedata             (mm_interconnect_3_vector_controller_master_0_slave_writedata), //                      .writedata
		.irq                         (irq_mapper_receiver4_irq)                                      //                   irq.irq
	);

	controller_vic_0 vic_0 (
		.clk_clk                        (clk_sys_clk),                                  //                      clk.clk
		.reset_reset                    (rst_controller_001_reset_out_reset),           //                    reset.reset
		.irq_input_irq                  (vic_0_irq_input_irq),                          //                irq_input.irq
		.csr_access_read                (mm_interconnect_2_vic_0_csr_access_read),      //               csr_access.read
		.csr_access_write               (mm_interconnect_2_vic_0_csr_access_write),     //                         .write
		.csr_access_address             (mm_interconnect_2_vic_0_csr_access_address),   //                         .address
		.csr_access_writedata           (mm_interconnect_2_vic_0_csr_access_writedata), //                         .writedata
		.csr_access_readdata            (mm_interconnect_2_vic_0_csr_access_readdata),  //                         .readdata
		.interrupt_controller_out_valid (vic_0_interrupt_controller_out_valid),         // interrupt_controller_out.valid
		.interrupt_controller_out_data  (vic_0_interrupt_controller_out_data)           //                         .data
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_0_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_0_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_0_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_0_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_0_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_0_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_0_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_0_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_0_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_0_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios_0_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios_0_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_0_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios_0_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios_0_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios_0_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios_0_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios_0_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios_0_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios_0_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios_0_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios_0_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios_0_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (nios_0_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (nios_0_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (nios_0_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (nios_0_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (nios_0_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (nios_0_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (nios_0_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (nios_0_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (nios_0_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (nios_0_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (nios_0_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (nios_0_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (nios_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_0_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	controller_nios_0_custom_instruction_master_comb_xconnect nios_0_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios_0_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios_0_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios_0_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios_0_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios_0_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios_0_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios_0_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios_0_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios_0_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios_0_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios_0_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios_0_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios_0_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios_0_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios_0_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios_0_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios_0_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios_0_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios_0_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios_0_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios_0_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_0_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_0_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_0_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_0_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_0_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_0_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_0_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios_0_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_clk       (),                                                                         // (terminated)
		.ci_master_clken     (),                                                                         // (terminated)
		.ci_master_reset_req (),                                                                         // (terminated)
		.ci_master_reset     (),                                                                         // (terminated)
		.ci_master_start     (),                                                                         // (terminated)
		.ci_master_done      (1'b0),                                                                     // (terminated)
		.ci_slave_clk        (1'b0),                                                                     // (terminated)
		.ci_slave_clken      (1'b0),                                                                     // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                     // (terminated)
		.ci_slave_reset      (1'b0),                                                                     // (terminated)
		.ci_slave_start      (1'b0),                                                                     // (terminated)
		.ci_slave_done       ()                                                                          // (terminated)
	);

	controller_nios_0_custom_instruction_master_multi_xconnect nios_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                      //           .ipending
		.ci_slave_estatus     (),                                                                      //           .estatus
		.ci_slave_clk         (nios_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios_0_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios_0_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios_0_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios_0_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios_0_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios_0_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_0_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_0_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_0_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_0_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios_0_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios_0_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_datab     (),                                                                          // (terminated)
		.ci_master_n         (),                                                                          // (terminated)
		.ci_master_readra    (),                                                                          // (terminated)
		.ci_master_readrb    (),                                                                          // (terminated)
		.ci_master_writerc   (),                                                                          // (terminated)
		.ci_master_a         (),                                                                          // (terminated)
		.ci_master_b         (),                                                                          // (terminated)
		.ci_master_c         (),                                                                          // (terminated)
		.ci_master_ipending  (),                                                                          // (terminated)
		.ci_master_estatus   (),                                                                          // (terminated)
		.ci_master_reset_req ()                                                                           // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios_0_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_datab),             //          .datab
		.ci_slave_result     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_result),            //          .result
		.ci_slave_n          (nios_0_custom_instruction_master_multi_xconnect_ci_master1_n),                 //          .n
		.ci_slave_readra     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_readra),            //          .readra
		.ci_slave_readrb     (nios_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),            //          .readrb
		.ci_slave_writerc    (nios_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),           //          .writerc
		.ci_slave_a          (nios_0_custom_instruction_master_multi_xconnect_ci_master1_a),                 //          .a
		.ci_slave_b          (nios_0_custom_instruction_master_multi_xconnect_ci_master1_b),                 //          .b
		.ci_slave_c          (nios_0_custom_instruction_master_multi_xconnect_ci_master1_c),                 //          .c
		.ci_slave_ipending   (nios_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),          //          .ipending
		.ci_slave_estatus    (nios_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),           //          .estatus
		.ci_slave_clk        (nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk),               //          .clk
		.ci_slave_clken      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),            //          .clk_en
		.ci_slave_reset_req  (nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),         //          .reset_req
		.ci_slave_reset      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_reset),             //          .reset
		.ci_slave_start      (nios_0_custom_instruction_master_multi_xconnect_ci_master1_start),             //          .start
		.ci_slave_done       (nios_0_custom_instruction_master_multi_xconnect_ci_master1_done),              //          .done
		.ci_master_dataa     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),     //          .datab
		.ci_master_result    (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_result),    //          .result
		.ci_master_n         (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_n),         //          .n
		.ci_master_clk       (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),       //          .clk
		.ci_master_clken     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),     //          .reset
		.ci_master_start     (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_start),     //          .start
		.ci_master_done      (nios_0_custom_instruction_master_multi_slave_translator1_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   ()                                                                              // (terminated)
	);

	controller_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                                (clk_sys_clk),                                                        //                                                              clk_0_clk.clk
		.spi_slave_to_avalon_mm_master_bridge_0_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // spi_slave_to_avalon_mm_master_bridge_0_clk_reset_reset_bridge_in_reset.reset
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address                 (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_address),       //                   spi_slave_to_avalon_mm_master_bridge_0_avalon_master.address
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest             (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_waitrequest),   //                                                                       .waitrequest
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable              (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_byteenable),    //                                                                       .byteenable
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read                    (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_read),          //                                                                       .read
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata                (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdata),      //                                                                       .readdata
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid           (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_readdatavalid), //                                                                       .readdatavalid
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write                   (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_write),         //                                                                       .write
		.spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata               (spi_slave_to_avalon_mm_master_bridge_0_avalon_master_writedata),     //                                                                       .writedata
		.data_ram_1_s2_address                                                        (mm_interconnect_0_data_ram_1_s2_address),                            //                                                          data_ram_1_s2.address
		.data_ram_1_s2_write                                                          (mm_interconnect_0_data_ram_1_s2_write),                              //                                                                       .write
		.data_ram_1_s2_readdata                                                       (mm_interconnect_0_data_ram_1_s2_readdata),                           //                                                                       .readdata
		.data_ram_1_s2_writedata                                                      (mm_interconnect_0_data_ram_1_s2_writedata),                          //                                                                       .writedata
		.data_ram_1_s2_byteenable                                                     (mm_interconnect_0_data_ram_1_s2_byteenable),                         //                                                                       .byteenable
		.data_ram_1_s2_chipselect                                                     (mm_interconnect_0_data_ram_1_s2_chipselect),                         //                                                                       .chipselect
		.data_ram_1_s2_clken                                                          (mm_interconnect_0_data_ram_1_s2_clken),                              //                                                                       .clken
		.mm_bridge_2_s0_address                                                       (mm_interconnect_0_mm_bridge_2_s0_address),                           //                                                         mm_bridge_2_s0.address
		.mm_bridge_2_s0_write                                                         (mm_interconnect_0_mm_bridge_2_s0_write),                             //                                                                       .write
		.mm_bridge_2_s0_read                                                          (mm_interconnect_0_mm_bridge_2_s0_read),                              //                                                                       .read
		.mm_bridge_2_s0_readdata                                                      (mm_interconnect_0_mm_bridge_2_s0_readdata),                          //                                                                       .readdata
		.mm_bridge_2_s0_writedata                                                     (mm_interconnect_0_mm_bridge_2_s0_writedata),                         //                                                                       .writedata
		.mm_bridge_2_s0_burstcount                                                    (mm_interconnect_0_mm_bridge_2_s0_burstcount),                        //                                                                       .burstcount
		.mm_bridge_2_s0_byteenable                                                    (mm_interconnect_0_mm_bridge_2_s0_byteenable),                        //                                                                       .byteenable
		.mm_bridge_2_s0_readdatavalid                                                 (mm_interconnect_0_mm_bridge_2_s0_readdatavalid),                     //                                                                       .readdatavalid
		.mm_bridge_2_s0_waitrequest                                                   (mm_interconnect_0_mm_bridge_2_s0_waitrequest),                       //                                                                       .waitrequest
		.mm_bridge_2_s0_debugaccess                                                   (mm_interconnect_0_mm_bridge_2_s0_debugaccess)                        //                                                                       .debugaccess
	);

	controller_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                        (clk_sys_clk),                                          //                                      clk_0_clk.clk
		.instruction_rom_0_reset1_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // instruction_rom_0_reset1_reset_bridge_in_reset.reset
		.mm_bridge_1_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                   //        mm_bridge_1_reset_reset_bridge_in_reset.reset
		.nios_0_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                   //             nios_0_reset_reset_bridge_in_reset.reset
		.nios_0_data_master_address                           (nios_0_data_master_address),                           //                             nios_0_data_master.address
		.nios_0_data_master_waitrequest                       (nios_0_data_master_waitrequest),                       //                                               .waitrequest
		.nios_0_data_master_byteenable                        (nios_0_data_master_byteenable),                        //                                               .byteenable
		.nios_0_data_master_read                              (nios_0_data_master_read),                              //                                               .read
		.nios_0_data_master_readdata                          (nios_0_data_master_readdata),                          //                                               .readdata
		.nios_0_data_master_write                             (nios_0_data_master_write),                             //                                               .write
		.nios_0_data_master_writedata                         (nios_0_data_master_writedata),                         //                                               .writedata
		.nios_0_data_master_debugaccess                       (nios_0_data_master_debugaccess),                       //                                               .debugaccess
		.nios_0_instruction_master_address                    (nios_0_instruction_master_address),                    //                      nios_0_instruction_master.address
		.nios_0_instruction_master_waitrequest                (nios_0_instruction_master_waitrequest),                //                                               .waitrequest
		.nios_0_instruction_master_read                       (nios_0_instruction_master_read),                       //                                               .read
		.nios_0_instruction_master_readdata                   (nios_0_instruction_master_readdata),                   //                                               .readdata
		.data_ram_0_s1_address                                (mm_interconnect_1_data_ram_0_s1_address),              //                                  data_ram_0_s1.address
		.data_ram_0_s1_write                                  (mm_interconnect_1_data_ram_0_s1_write),                //                                               .write
		.data_ram_0_s1_readdata                               (mm_interconnect_1_data_ram_0_s1_readdata),             //                                               .readdata
		.data_ram_0_s1_writedata                              (mm_interconnect_1_data_ram_0_s1_writedata),            //                                               .writedata
		.data_ram_0_s1_byteenable                             (mm_interconnect_1_data_ram_0_s1_byteenable),           //                                               .byteenable
		.data_ram_0_s1_chipselect                             (mm_interconnect_1_data_ram_0_s1_chipselect),           //                                               .chipselect
		.data_ram_0_s1_clken                                  (mm_interconnect_1_data_ram_0_s1_clken),                //                                               .clken
		.data_ram_1_s1_address                                (mm_interconnect_1_data_ram_1_s1_address),              //                                  data_ram_1_s1.address
		.data_ram_1_s1_write                                  (mm_interconnect_1_data_ram_1_s1_write),                //                                               .write
		.data_ram_1_s1_readdata                               (mm_interconnect_1_data_ram_1_s1_readdata),             //                                               .readdata
		.data_ram_1_s1_writedata                              (mm_interconnect_1_data_ram_1_s1_writedata),            //                                               .writedata
		.data_ram_1_s1_byteenable                             (mm_interconnect_1_data_ram_1_s1_byteenable),           //                                               .byteenable
		.data_ram_1_s1_chipselect                             (mm_interconnect_1_data_ram_1_s1_chipselect),           //                                               .chipselect
		.data_ram_1_s1_clken                                  (mm_interconnect_1_data_ram_1_s1_clken),                //                                               .clken
		.instruction_rom_0_s1_address                         (mm_interconnect_1_instruction_rom_0_s1_address),       //                           instruction_rom_0_s1.address
		.instruction_rom_0_s1_write                           (mm_interconnect_1_instruction_rom_0_s1_write),         //                                               .write
		.instruction_rom_0_s1_readdata                        (mm_interconnect_1_instruction_rom_0_s1_readdata),      //                                               .readdata
		.instruction_rom_0_s1_writedata                       (mm_interconnect_1_instruction_rom_0_s1_writedata),     //                                               .writedata
		.instruction_rom_0_s1_byteenable                      (mm_interconnect_1_instruction_rom_0_s1_byteenable),    //                                               .byteenable
		.instruction_rom_0_s1_chipselect                      (mm_interconnect_1_instruction_rom_0_s1_chipselect),    //                                               .chipselect
		.instruction_rom_0_s1_clken                           (mm_interconnect_1_instruction_rom_0_s1_clken),         //                                               .clken
		.mm_bridge_0_s0_address                               (mm_interconnect_1_mm_bridge_0_s0_address),             //                                 mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                 (mm_interconnect_1_mm_bridge_0_s0_write),               //                                               .write
		.mm_bridge_0_s0_read                                  (mm_interconnect_1_mm_bridge_0_s0_read),                //                                               .read
		.mm_bridge_0_s0_readdata                              (mm_interconnect_1_mm_bridge_0_s0_readdata),            //                                               .readdata
		.mm_bridge_0_s0_writedata                             (mm_interconnect_1_mm_bridge_0_s0_writedata),           //                                               .writedata
		.mm_bridge_0_s0_burstcount                            (mm_interconnect_1_mm_bridge_0_s0_burstcount),          //                                               .burstcount
		.mm_bridge_0_s0_byteenable                            (mm_interconnect_1_mm_bridge_0_s0_byteenable),          //                                               .byteenable
		.mm_bridge_0_s0_readdatavalid                         (mm_interconnect_1_mm_bridge_0_s0_readdatavalid),       //                                               .readdatavalid
		.mm_bridge_0_s0_waitrequest                           (mm_interconnect_1_mm_bridge_0_s0_waitrequest),         //                                               .waitrequest
		.mm_bridge_0_s0_debugaccess                           (mm_interconnect_1_mm_bridge_0_s0_debugaccess),         //                                               .debugaccess
		.mm_bridge_1_s0_address                               (mm_interconnect_1_mm_bridge_1_s0_address),             //                                 mm_bridge_1_s0.address
		.mm_bridge_1_s0_write                                 (mm_interconnect_1_mm_bridge_1_s0_write),               //                                               .write
		.mm_bridge_1_s0_read                                  (mm_interconnect_1_mm_bridge_1_s0_read),                //                                               .read
		.mm_bridge_1_s0_readdata                              (mm_interconnect_1_mm_bridge_1_s0_readdata),            //                                               .readdata
		.mm_bridge_1_s0_writedata                             (mm_interconnect_1_mm_bridge_1_s0_writedata),           //                                               .writedata
		.mm_bridge_1_s0_burstcount                            (mm_interconnect_1_mm_bridge_1_s0_burstcount),          //                                               .burstcount
		.mm_bridge_1_s0_byteenable                            (mm_interconnect_1_mm_bridge_1_s0_byteenable),          //                                               .byteenable
		.mm_bridge_1_s0_readdatavalid                         (mm_interconnect_1_mm_bridge_1_s0_readdatavalid),       //                                               .readdatavalid
		.mm_bridge_1_s0_waitrequest                           (mm_interconnect_1_mm_bridge_1_s0_waitrequest),         //                                               .waitrequest
		.mm_bridge_1_s0_debugaccess                           (mm_interconnect_1_mm_bridge_1_s0_debugaccess),         //                                               .debugaccess
		.nios_0_debug_mem_slave_address                       (mm_interconnect_1_nios_0_debug_mem_slave_address),     //                         nios_0_debug_mem_slave.address
		.nios_0_debug_mem_slave_write                         (mm_interconnect_1_nios_0_debug_mem_slave_write),       //                                               .write
		.nios_0_debug_mem_slave_read                          (mm_interconnect_1_nios_0_debug_mem_slave_read),        //                                               .read
		.nios_0_debug_mem_slave_readdata                      (mm_interconnect_1_nios_0_debug_mem_slave_readdata),    //                                               .readdata
		.nios_0_debug_mem_slave_writedata                     (mm_interconnect_1_nios_0_debug_mem_slave_writedata),   //                                               .writedata
		.nios_0_debug_mem_slave_byteenable                    (mm_interconnect_1_nios_0_debug_mem_slave_byteenable),  //                                               .byteenable
		.nios_0_debug_mem_slave_waitrequest                   (mm_interconnect_1_nios_0_debug_mem_slave_waitrequest), //                                               .waitrequest
		.nios_0_debug_mem_slave_debugaccess                   (mm_interconnect_1_nios_0_debug_mem_slave_debugaccess)  //                                               .debugaccess
	);

	controller_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                           (clk_sys_clk),                                                         //                                         clk_0_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset           (rst_controller_003_reset_out_reset),                                  //           mm_bridge_0_reset_reset_bridge_in_reset.reset
		.performance_counter_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                  // performance_counter_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                                  (mm_bridge_0_m0_address),                                              //                                    mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                              (mm_bridge_0_m0_waitrequest),                                          //                                                  .waitrequest
		.mm_bridge_0_m0_burstcount                               (mm_bridge_0_m0_burstcount),                                           //                                                  .burstcount
		.mm_bridge_0_m0_byteenable                               (mm_bridge_0_m0_byteenable),                                           //                                                  .byteenable
		.mm_bridge_0_m0_read                                     (mm_bridge_0_m0_read),                                                 //                                                  .read
		.mm_bridge_0_m0_readdata                                 (mm_bridge_0_m0_readdata),                                             //                                                  .readdata
		.mm_bridge_0_m0_readdatavalid                            (mm_bridge_0_m0_readdatavalid),                                        //                                                  .readdatavalid
		.mm_bridge_0_m0_write                                    (mm_bridge_0_m0_write),                                                //                                                  .write
		.mm_bridge_0_m0_writedata                                (mm_bridge_0_m0_writedata),                                            //                                                  .writedata
		.mm_bridge_0_m0_debugaccess                              (mm_bridge_0_m0_debugaccess),                                          //                                                  .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address                   (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_address),             //                     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                     (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_write),               //                                                  .write
		.jtag_uart_0_avalon_jtag_slave_read                      (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_read),                //                                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata                  (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_readdata),            //                                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                 (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_writedata),           //                                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest               (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_waitrequest),         //                                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                (mm_interconnect_2_jtag_uart_0_avalon_jtag_slave_chipselect),          //                                                  .chipselect
		.msgdma_0_csr_address                                    (mm_interconnect_2_msgdma_0_csr_address),                              //                                      msgdma_0_csr.address
		.msgdma_0_csr_write                                      (mm_interconnect_2_msgdma_0_csr_write),                                //                                                  .write
		.msgdma_0_csr_read                                       (mm_interconnect_2_msgdma_0_csr_read),                                 //                                                  .read
		.msgdma_0_csr_readdata                                   (mm_interconnect_2_msgdma_0_csr_readdata),                             //                                                  .readdata
		.msgdma_0_csr_writedata                                  (mm_interconnect_2_msgdma_0_csr_writedata),                            //                                                  .writedata
		.msgdma_0_csr_byteenable                                 (mm_interconnect_2_msgdma_0_csr_byteenable),                           //                                                  .byteenable
		.msgdma_0_descriptor_slave_write                         (mm_interconnect_2_msgdma_0_descriptor_slave_write),                   //                         msgdma_0_descriptor_slave.write
		.msgdma_0_descriptor_slave_writedata                     (mm_interconnect_2_msgdma_0_descriptor_slave_writedata),               //                                                  .writedata
		.msgdma_0_descriptor_slave_byteenable                    (mm_interconnect_2_msgdma_0_descriptor_slave_byteenable),              //                                                  .byteenable
		.msgdma_0_descriptor_slave_waitrequest                   (mm_interconnect_2_msgdma_0_descriptor_slave_waitrequest),             //                                                  .waitrequest
		.performance_counter_0_control_slave_address             (mm_interconnect_2_performance_counter_0_control_slave_address),       //               performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write               (mm_interconnect_2_performance_counter_0_control_slave_write),         //                                                  .write
		.performance_counter_0_control_slave_readdata            (mm_interconnect_2_performance_counter_0_control_slave_readdata),      //                                                  .readdata
		.performance_counter_0_control_slave_writedata           (mm_interconnect_2_performance_counter_0_control_slave_writedata),     //                                                  .writedata
		.performance_counter_0_control_slave_begintransfer       (mm_interconnect_2_performance_counter_0_control_slave_begintransfer), //                                                  .begintransfer
		.sysid_qsys_0_control_slave_address                      (mm_interconnect_2_sysid_qsys_0_control_slave_address),                //                        sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                     (mm_interconnect_2_sysid_qsys_0_control_slave_readdata),               //                                                  .readdata
		.timer_0_s1_address                                      (mm_interconnect_2_timer_0_s1_address),                                //                                        timer_0_s1.address
		.timer_0_s1_write                                        (mm_interconnect_2_timer_0_s1_write),                                  //                                                  .write
		.timer_0_s1_readdata                                     (mm_interconnect_2_timer_0_s1_readdata),                               //                                                  .readdata
		.timer_0_s1_writedata                                    (mm_interconnect_2_timer_0_s1_writedata),                              //                                                  .writedata
		.timer_0_s1_chipselect                                   (mm_interconnect_2_timer_0_s1_chipselect),                             //                                                  .chipselect
		.vic_0_csr_access_address                                (mm_interconnect_2_vic_0_csr_access_address),                          //                                  vic_0_csr_access.address
		.vic_0_csr_access_write                                  (mm_interconnect_2_vic_0_csr_access_write),                            //                                                  .write
		.vic_0_csr_access_read                                   (mm_interconnect_2_vic_0_csr_access_read),                             //                                                  .read
		.vic_0_csr_access_readdata                               (mm_interconnect_2_vic_0_csr_access_readdata),                         //                                                  .readdata
		.vic_0_csr_access_writedata                              (mm_interconnect_2_vic_0_csr_access_writedata)                         //                                                  .writedata
	);

	controller_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                        (clk_sys_clk),                                                  //                                      clk_0_clk.clk
		.mm_bridge_1_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                           //        mm_bridge_1_reset_reset_bridge_in_reset.reset
		.motor_controller_5_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // motor_controller_5_reset_reset_bridge_in_reset.reset
		.mm_bridge_1_m0_address                               (mm_bridge_1_m0_address),                                       //                                 mm_bridge_1_m0.address
		.mm_bridge_1_m0_waitrequest                           (mm_bridge_1_m0_waitrequest),                                   //                                               .waitrequest
		.mm_bridge_1_m0_burstcount                            (mm_bridge_1_m0_burstcount),                                    //                                               .burstcount
		.mm_bridge_1_m0_byteenable                            (mm_bridge_1_m0_byteenable),                                    //                                               .byteenable
		.mm_bridge_1_m0_read                                  (mm_bridge_1_m0_read),                                          //                                               .read
		.mm_bridge_1_m0_readdata                              (mm_bridge_1_m0_readdata),                                      //                                               .readdata
		.mm_bridge_1_m0_readdatavalid                         (mm_bridge_1_m0_readdatavalid),                                 //                                               .readdatavalid
		.mm_bridge_1_m0_write                                 (mm_bridge_1_m0_write),                                         //                                               .write
		.mm_bridge_1_m0_writedata                             (mm_bridge_1_m0_writedata),                                     //                                               .writedata
		.mm_bridge_1_m0_debugaccess                           (mm_bridge_1_m0_debugaccess),                                   //                                               .debugaccess
		.i2c_master_0_slave_address                           (mm_interconnect_3_i2c_master_0_slave_address),                 //                             i2c_master_0_slave.address
		.i2c_master_0_slave_write                             (mm_interconnect_3_i2c_master_0_slave_write),                   //                                               .write
		.i2c_master_0_slave_read                              (mm_interconnect_3_i2c_master_0_slave_read),                    //                                               .read
		.i2c_master_0_slave_readdata                          (mm_interconnect_3_i2c_master_0_slave_readdata),                //                                               .readdata
		.i2c_master_0_slave_writedata                         (mm_interconnect_3_i2c_master_0_slave_writedata),               //                                               .writedata
		.imu_spim_slave_address                               (mm_interconnect_3_imu_spim_slave_address),                     //                                 imu_spim_slave.address
		.imu_spim_slave_write                                 (mm_interconnect_3_imu_spim_slave_write),                       //                                               .write
		.imu_spim_slave_read                                  (mm_interconnect_3_imu_spim_slave_read),                        //                                               .read
		.imu_spim_slave_readdata                              (mm_interconnect_3_imu_spim_slave_readdata),                    //                                               .readdata
		.imu_spim_slave_writedata                             (mm_interconnect_3_imu_spim_slave_writedata),                   //                                               .writedata
		.motor_controller_5_slave_address                     (mm_interconnect_3_motor_controller_5_slave_address),           //                       motor_controller_5_slave.address
		.motor_controller_5_slave_write                       (mm_interconnect_3_motor_controller_5_slave_write),             //                                               .write
		.motor_controller_5_slave_read                        (mm_interconnect_3_motor_controller_5_slave_read),              //                                               .read
		.motor_controller_5_slave_readdata                    (mm_interconnect_3_motor_controller_5_slave_readdata),          //                                               .readdata
		.motor_controller_5_slave_writedata                   (mm_interconnect_3_motor_controller_5_slave_writedata),         //                                               .writedata
		.pio_0_s1_address                                     (mm_interconnect_3_pio_0_s1_address),                           //                                       pio_0_s1.address
		.pio_0_s1_write                                       (mm_interconnect_3_pio_0_s1_write),                             //                                               .write
		.pio_0_s1_readdata                                    (mm_interconnect_3_pio_0_s1_readdata),                          //                                               .readdata
		.pio_0_s1_writedata                                   (mm_interconnect_3_pio_0_s1_writedata),                         //                                               .writedata
		.pio_0_s1_chipselect                                  (mm_interconnect_3_pio_0_s1_chipselect),                        //                                               .chipselect
		.pio_1_s1_address                                     (mm_interconnect_3_pio_1_s1_address),                           //                                       pio_1_s1.address
		.pio_1_s1_write                                       (mm_interconnect_3_pio_1_s1_write),                             //                                               .write
		.pio_1_s1_readdata                                    (mm_interconnect_3_pio_1_s1_readdata),                          //                                               .readdata
		.pio_1_s1_writedata                                   (mm_interconnect_3_pio_1_s1_writedata),                         //                                               .writedata
		.pio_1_s1_chipselect                                  (mm_interconnect_3_pio_1_s1_chipselect),                        //                                               .chipselect
		.pio_2_s1_address                                     (mm_interconnect_3_pio_2_s1_address),                           //                                       pio_2_s1.address
		.pio_2_s1_write                                       (mm_interconnect_3_pio_2_s1_write),                             //                                               .write
		.pio_2_s1_readdata                                    (mm_interconnect_3_pio_2_s1_readdata),                          //                                               .readdata
		.pio_2_s1_writedata                                   (mm_interconnect_3_pio_2_s1_writedata),                         //                                               .writedata
		.pio_2_s1_chipselect                                  (mm_interconnect_3_pio_2_s1_chipselect),                        //                                               .chipselect
		.spim_0_spi_control_port_address                      (mm_interconnect_3_spim_0_spi_control_port_address),            //                        spim_0_spi_control_port.address
		.spim_0_spi_control_port_write                        (mm_interconnect_3_spim_0_spi_control_port_write),              //                                               .write
		.spim_0_spi_control_port_read                         (mm_interconnect_3_spim_0_spi_control_port_read),               //                                               .read
		.spim_0_spi_control_port_readdata                     (mm_interconnect_3_spim_0_spi_control_port_readdata),           //                                               .readdata
		.spim_0_spi_control_port_writedata                    (mm_interconnect_3_spim_0_spi_control_port_writedata),          //                                               .writedata
		.spim_0_spi_control_port_chipselect                   (mm_interconnect_3_spim_0_spi_control_port_chipselect),         //                                               .chipselect
		.vector_controller_master_0_slave_address             (mm_interconnect_3_vector_controller_master_0_slave_address),   //               vector_controller_master_0_slave.address
		.vector_controller_master_0_slave_write               (mm_interconnect_3_vector_controller_master_0_slave_write),     //                                               .write
		.vector_controller_master_0_slave_read                (mm_interconnect_3_vector_controller_master_0_slave_read),      //                                               .read
		.vector_controller_master_0_slave_readdata            (mm_interconnect_3_vector_controller_master_0_slave_readdata),  //                                               .readdata
		.vector_controller_master_0_slave_writedata           (mm_interconnect_3_vector_controller_master_0_slave_writedata)  //                                               .writedata
	);

	controller_mm_interconnect_4 mm_interconnect_4 (
		.clk_0_clk_clk                                 (clk_sys_clk),                                       //                               clk_0_clk.clk
		.mm_bridge_2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // mm_bridge_2_reset_reset_bridge_in_reset.reset
		.msgdma_0_reset_n_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                //  msgdma_0_reset_n_reset_bridge_in_reset.reset
		.mm_bridge_2_m0_address                        (mm_bridge_2_m0_address),                            //                          mm_bridge_2_m0.address
		.mm_bridge_2_m0_waitrequest                    (mm_bridge_2_m0_waitrequest),                        //                                        .waitrequest
		.mm_bridge_2_m0_burstcount                     (mm_bridge_2_m0_burstcount),                         //                                        .burstcount
		.mm_bridge_2_m0_byteenable                     (mm_bridge_2_m0_byteenable),                         //                                        .byteenable
		.mm_bridge_2_m0_read                           (mm_bridge_2_m0_read),                               //                                        .read
		.mm_bridge_2_m0_readdata                       (mm_bridge_2_m0_readdata),                           //                                        .readdata
		.mm_bridge_2_m0_readdatavalid                  (mm_bridge_2_m0_readdatavalid),                      //                                        .readdatavalid
		.mm_bridge_2_m0_write                          (mm_bridge_2_m0_write),                              //                                        .write
		.mm_bridge_2_m0_writedata                      (mm_bridge_2_m0_writedata),                          //                                        .writedata
		.mm_bridge_2_m0_debugaccess                    (mm_bridge_2_m0_debugaccess),                        //                                        .debugaccess
		.msgdma_0_mm_read_address                      (msgdma_0_mm_read_address),                          //                        msgdma_0_mm_read.address
		.msgdma_0_mm_read_waitrequest                  (msgdma_0_mm_read_waitrequest),                      //                                        .waitrequest
		.msgdma_0_mm_read_read                         (msgdma_0_mm_read_read),                             //                                        .read
		.msgdma_0_mm_read_readdata                     (msgdma_0_mm_read_readdata),                         //                                        .readdata
		.msgdma_0_mm_read_readdatavalid                (msgdma_0_mm_read_readdatavalid),                    //                                        .readdatavalid
		.data_ram_0_s2_address                         (mm_interconnect_4_data_ram_0_s2_address),           //                           data_ram_0_s2.address
		.data_ram_0_s2_write                           (mm_interconnect_4_data_ram_0_s2_write),             //                                        .write
		.data_ram_0_s2_readdata                        (mm_interconnect_4_data_ram_0_s2_readdata),          //                                        .readdata
		.data_ram_0_s2_writedata                       (mm_interconnect_4_data_ram_0_s2_writedata),         //                                        .writedata
		.data_ram_0_s2_byteenable                      (mm_interconnect_4_data_ram_0_s2_byteenable),        //                                        .byteenable
		.data_ram_0_s2_chipselect                      (mm_interconnect_4_data_ram_0_s2_chipselect),        //                                        .chipselect
		.data_ram_0_s2_clken                           (mm_interconnect_4_data_ram_0_s2_clken),             //                                        .clken
		.instruction_rom_0_s2_address                  (mm_interconnect_4_instruction_rom_0_s2_address),    //                    instruction_rom_0_s2.address
		.instruction_rom_0_s2_write                    (mm_interconnect_4_instruction_rom_0_s2_write),      //                                        .write
		.instruction_rom_0_s2_readdata                 (mm_interconnect_4_instruction_rom_0_s2_readdata),   //                                        .readdata
		.instruction_rom_0_s2_writedata                (mm_interconnect_4_instruction_rom_0_s2_writedata),  //                                        .writedata
		.instruction_rom_0_s2_byteenable               (mm_interconnect_4_instruction_rom_0_s2_byteenable), //                                        .byteenable
		.instruction_rom_0_s2_chipselect               (mm_interconnect_4_instruction_rom_0_s2_chipselect), //                                        .chipselect
		.instruction_rom_0_s2_clken                    (mm_interconnect_4_instruction_rom_0_s2_clken)       //                                        .clken
	);

	controller_irq_mapper irq_mapper (
		.clk           (clk_sys_clk),                        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),           // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),           // receiver8.irq
		.sender_irq    (vic_0_irq_input_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_sys_reset_n),                 // reset_in0.reset
		.clk            (clk_sys_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_sys_reset_n),                 // reset_in0.reset
		.reset_in1      (nios_0_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (reset_controller_0_reset_out_reset), // reset_in2.reset
		.clk            (clk_sys_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_100mhz_reset_n),              // reset_in0.reset
		.clk            (clk_100mhz_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_sys_reset_n),                     // reset_in0.reset
		.reset_in1      (reset_controller_0_reset_out_reset),     // reset_in1.reset
		.clk            (clk_sys_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_sys_reset_n),                 // reset_in0.reset
		.reset_in1      (nios_0_debug_reset_request_reset),   // reset_in1.reset
		.reset_in2      (reset_controller_0_reset_out_reset), // reset_in2.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
