// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 14:37:35 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
chCtv9yLoUaSv6+wD+pSyubsXklt96maOqwIbzT0sXbR9xD7OD0MSy/JSXCnWCYq
XR0OXGS/abG1mqIzOJAURbOUxfBuhTPEdFpzBj412NATSPelg6Bz8IEUh3vMFtbh
HmTTUMHU0svRZpv/weUn06O1WTzZsvDjtHbWa3WxrEQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
NsM27Wi4UGBNQAXmgtc2Zx3BytEpxqAzuPJk9/3zHlBqmrS7gWCsXgZjAjaSqpmC
IDG5cb1e+LVWCeax1rF0dmbhdru+7rLnFxdQ433dC9/++KvD3NDlIK7gSq3fi3Zh
9eNzh/Lc4Q5VUr2xIwTgBXE6ZywFRqULlCBqDUMXt3uwfTgUBl7x7Ord/EnjUDc1
UdV60Hy8H+AXg5U1k/QdCyPJuVcmzgvU/mvxapg5XFJ8GgSKB06U4FsH/pjXvfbM
1BusefU9E9MvFq8CqM8OeOvyh6TATfZEJlKg7HO3Glbl8QdSBeC5zSoHI/ACaxVW
lJBsp5vWqSM0hMJI4q7iKOegIyAIXV3/mwq/rKdfqhhfTGyA3/D7MzWa0+nbcr76
aurAcU2Mw0uQ42pDVJoETflJ6dy0CwCK9CZaE2s3u/HVvuEyDH1QWisJqFHPm0kh
TIzhmjCUdqOIiKuJDfE0zgqgq7+bDMRVzdFAJqlbmCUDW3YwTu8rKii2ZsxKUhLs
CZNc37CQYVEP7a+PPKi4SVFSV2NAOfD/C65va4Y28NwY9Kf+048PKOn4cYxuL1xv
5KS2iR+gV7z16fKAv0Hr8RY5eE3LjpJ5xahr6ybK/PzV+1dcr7ddi37HAwlLx58i
akvKGCYILeZDsmiUc5owRke8aJDeJ2KyEJh0uTG/Uj7DHClzkjrEbvZ0QbgY1KYa
KqMznHlzttnWrNwIOe7znW+/9RM3UXNQKxUyXaI0Fx1g5RNwtXkHXRrGZcPDYU1f
pw7vFU/+CzlhuffTopDMfW/Xo5L238QPjtJXXc9f4aqWVwR8Wwt6nlb20zw1jsXh
6FcdEBLCD6o54eoxqxsw0B7x49lFltcb0CajY+ufB0rC+cVtDXo363pPvW0yXe+C
ibZbZ+SYhVyOUPeaoGkkeBITykvolIhX3o4V7jMgCzAp9mmaiN/DiEqdZcbw4CdI
TwsD3P/CvAEuEYptOl+CqkKtnFnjc0jTXbFCA6IgqsVIJTdghk+HaEdV0fN9QyaM
bLVc19KPAnrodG8hrtp2Cs0kh4HGKWh8oX1c8zon3CaXsB52kHV4pvpfNv2SA09o
3OzYGhNXkBbIfFxc6MI9CZoaU5sFI9vkua13BQxIQ/BWwW3CIAsotjDkrEx5bUB1
vcoLV2iuEnD893XcqVMSXzvQ5f5PNsvA+we7mCvtf6D6Y2FeRH+vmCFZ3WCBTIR3
0Q9hi+73h/t3h0Alx07lOTNddWZCwpMi6jaew+6k0WtYxUjWu+9WUoKsjv6GSgIj
Y4D1t3/Btq4b9ZfNRP//2p/YwuknAO1MehxI6StxiUsGPsnRfwVEgUK/nRZh5Z8D
9uz1slzMxG9SoaQnODpuo4JUIRQ168U+swTCLtRnzuhi8oQRXBFF0goGWZFVDg7V
Ap9DsL5geFKzGBFoiqUZuyLaT25cOZh9ccC0gVVIkvn/cYNV7RrV+6m4db/SW/WV
QGJPPbOhP6dZ9mAV2UWw9EauL43zZR/F+kNrBO0waHhsOUx/tFcyuLKChdxds5mr
BGYoDEIWY91LrdoQa13w85TzzKXRagdiZGlpzr9vtp42XZnl22xmWA3vqPmISRvH
CbZ5sb02Tez34udsizxLNNU5ZMqduuxmb4iKUVGzQsUtC0zU1id0ZZEonPkGyc5R
PciXx/6BnXhvoN82096vs4v7ZnWKnVQ6zwhYJKnGpiFns3xR403VVMBRB55js8w2
QV6ME8i9IzZZVrAEvY9CTQG4Eh0HJlgCQ239eU4+eaArrjS/NJet8ftbAdybRpVB
JXaXDy0lGMd/xDDyHoI0/8MucgfvWgNcEadyisG86Efqp4cfGeU2jYXHy+rEM14h
zMf8NkhESNXG7hMerivnEqIr+j6LjEZxLQ/NjjJc4tCVCMX4L+dqwzph48s55Q9b
/K1shsI85AgrgcGYvLYOcc1mismYzItV5Y0TiEYf+Udr/0Cq+H19bpvP36NFwHTr
TxN1Mw66MUvlwNdV3BCGE7QsFsRchUlMVGn5gwBH5ghSmtCsNyjfMYlAi7BZbij5
6UjnpPt8R23dlsWP+D+DqkGr8EGNDifQLAcVbYRYTt8A0inTMrKeOL/PIrQ1YKBg
l8eqb9iS0d6siiapfOrq/2wZEPyJJ0gHwUqrDVqchRYHcyHlT03Gk0why0oCFmVS
uA3PUChpaeqd/blulTlQoZKrL72k7w1i+gI3gZLbL2zvrrXF5ihpUOyiLbIT9rz8
LH/y4G4/CuenZ3Kygu5jXhamGSDJ6oskTPtTgETeexmQZVI/Gz75fOVZ9dwNJP24
tkD/2OGb4ufRV/w0hpZke4rTmK2EED1R8YkSOkpRVH7oBkEI7wA8Arx1KOvauYs3
mqDPkuacQEzF6UTEEH8BiTAZ069n1J4Kwlm8lLs3D2mLFSaFRkxFuEP41z4vXFk1
PomBf8H6llXdcIazJ5M8vglR8lNG7m642AaFicLnMlOM87hQTH+nXxnaGDXHIlPM
Zq8df1lXwTucZ2polCNI+8vSge9LT7FzkQXewahzrNZCYekTwSd1BfdlkFqcVA8L
egQYpmrzK8Jm+jyOdr523PmcRgiihwIJB+MdYBoHlsph1TPcu2VvsUI02MSUNHlT
dblFBX+2lbuPczWNrj47Jghm132JcEk5VU5f3iLZpcy7yYuWKN2jOAxkOy2FW80v
k/VClEq2mDRnQLcE7vOdTHGckYlwwmolpUCI13FnffTp09vg+/yDa01T1h+BAUfG
tbS0umJBMOChwZAFUH50HuFlPPH4SD0kRfN7S5vFqrhy9qSEfqjIJZUJxpNb4EDL
8RhKfLZKxEESURF12h5nM7K3PK3LGCCYSDxku0VdO5DdKsti4Rbx0JFVrhE1owzQ
9YTeUVHa0rFSbU+gbSzIzUmIcLRk8l9N5G8jaTrANT9SnelL1xz6gVw3KmFYXhp+
3O6c6jV5L20OHMnHMrF8IozByVMDziPmMJcwezK5/Xcws8Tjl+xHlEUmsnpYB/bp
AzwRunuNSxBi5kwBZEdDoOzisQabsrf9loxFg8HKgBRW/KyBSA+Pqe4nHie0Q6Pv
e0F3F1Lhhcv6p3JpfcmIRVpJRbp/CAKy0oNF7DQ66jEh8C/splWsVv/2wdOUzkl5
3lkepNowdqtR0TOnx56fzhyANTi26Ike/H++LaHq96/KUFHQ2b2MkDJFfMwGoog/
0yzeldF3e/vPKv3eA8CbPo+NXBFR7TyuEzRa4iTzEiTSPZwKlbZmf660EJxECcuF
h5QiqGsAhsz82RrPMDfetZe5tJ3QtQ7vlo2yDuONXDLq0qKznU/mpIjk2uCFZs/I
nI6MDDAFIrrUPuQIqkCiMq1mFQkAx55AAZG90Q0uTxC/0VSt0qufAmxdOIDbWix2
a4gmGav+UgAvtA6PdB5crQflkbmxEIJB7z0kg8k5KYB57h72AlB7xHtaZtLyMGDr
ctPNIfm0h69xVkZbSI6X53U6TNd81Xo6p37zXmtxlfsLpExovdFLoBG0Wb7FO0m9
m4wGR5e8FBsSSQZFlcf3X9GcGt1wBPiK3faYbhHk30R1Kef0DXVQy6RuXLgEpTmq
ETmNmo47nhZjN7vNo1hjM33XrAZQT4Ucznljc3LA+7lws/210Bcu3Bo8KXC1HwrK
3Z7vjv6QjxVeHIperg9YPW6pgxK3l9QlKcfU00ywt7AnMUGGw+vi2ZRIVsom1eEW
e/M7ay7CWDKqyn57JGyo5seEqT2En4FVlD85kY2mGS28YYDHnpkibiofVk2EsPKB
cCFXE6FaV4dzg1EP3vZYWhfEoyhCK11oYBXwnsor43lDZ9HPQLgLsZFdYHLBik9r
8YliJ2fCdNz1gD0KB/ZB3egQIVmUrSUHqj0ZpjlXf5BuL6oW1GWKeAJlKJd38LEB
SyvPigOTrv/MU/L9ztxj3ti3j423nRMVNW4O5bl5cSDeMhvmFQ9PEUzbgWSoyUOr
5gem/MjOXJseKVpZH+dknmTrOnGt6Xvk1XPTqwJ6WSv0jBIQcWI96u2B/6qy9jJm
Fm/jqeReVbjAyYevszsmOyVrmagneDdiPNLVPK6Vn5DOYpUooV3BmXHpWX+Ur1Wb
hThkJFedzbs1sCrlwyzHrSit0x/7kmCLpgV6dXCHQpujg674Inuh+ZlePF3ttiaE
D68KPC/tNG8EAzXQb8CGYvvKRe3nW7wJoYx1MCS4GK1rmlPEHW9AjXKxYM/riXVD
EcDVYtmIO3FYxcZm05uAmDKgc1mLud37e2D2FcRIStT8BYiKo2suCdKk14U34C5T
kSdfTEMX3o8EAIwfrijFt4Nk5dDNuwUowLaJHWzHxuxSRDBi94DG1dST4d89LF2e
P7V8oCeB21W1tAkrU6phjfUcgqmLxEWCPxg6qM5zaDxFuqjsaPS9kRXMSD6OPZj/
E3SZtF2h9mzFj1N0aI4ocaMaBK7ARlmmkk/FPRRZj/Jg2GnwY1MRArtgLinnCA9z
s0DvJ1rVqKOyrlIRlgUtad4r6bIzvknme3jtFw+h+xo29tW2UWDARoW7IoE8CPvi
FtlTCtarDKfJlSS7TXaniybMqaq41bsRAFzbkkxGkOMHjYIDyDKs36DZ9UBoqVKq
+3ejnpf8gZgxzTk+1G7homQWKCCAXuimKyTXwSd4mvl/SIGx4CELaOzu+z2arIbY
UmE9u4HO8WKMbhVgyNwL8AhkggOeV14/rHAIxh8XaAsjRIz16dqw2U+i5EW18iLu
Ce3/qgbnniMwVOc6599TG9/BtCDOSNU7U1N/iZYldQw5YSyTm9EIe+lgRucjCHhZ
85mPX7bQVMg5i/BI88wGEdzQF4eHJaLV0d4XEpvhYamLQFpfzSsU7Txpp/65TmKx
vdUCQtyFJPBYtDePj28Z/RRUPDwIbr/MIMzE4dN7J2eHUUgAay+NEHiyD0WHPRO8
9JWgoQ9lcn9UnsSqaXSb4FL9z9MkdIsy6l/g3WuTcusmdX6fSrqhfFdpGw46S1hz
y8gxFAPvCF8I9RV8ghakDYb7k+Lr9IT65+HA0aDWLgnmL0xVKK0byPkbYGyFVgzX
E3/rZSbpYLPdzA/Wbro6ufWHIHaw7KGqDiPGOZQ4v6VsyjQ4kaFfsVYZTl6kgVlb
vRwFDaIV96xjbsMR0Y6Olxg6t7i4U4N6vNrlKa4LAjd6JSznl54tqBgcmZdnIllc
clL9jMhW0nAF+4SfOcxyPDZKQ5i8BqSgD0H3kFdRhQ5qTGsIJwDJgmrgBcz0+ncw
A7jaSOMSjGM6CG0RQQTWhDjKnPDdLF4uo5LpQA1XwbkKDbFXcHFoUq1eu+DLKEp0
jZE1L9yAdrgK7utx8ivtdORj3FofCGckIAuhck1rpLwQOoRB8IgFak9uKJtZOCzv
xKfETVL+GaVa431Ur2dmJBj5F6cwM9rBhhj0BE/T0wmsE05RxJ0bDxa36/usT1in
sLrp5DIB8I3HxExOx5oN7koSMWm5cY8DyEtTFEg+7E+HR9IutTF8la8KUrd/u+ZX
r6yttXVsKycbhgZaDXjoWdik+10jZMz8vZ48E3edpkfILKWgDSSFRlxQorU7/iUK
QezJBYcBe+uy5c3B5xSlz0TSLXnlcrjtNA6Nl9sQp59sWA/cAY3b9z8A4sjVfaKL
PlR8VaXcF+nJeRMomkpKPi+gjGMMjA8ZfLivCdK8lPSxPbMeqeYFPi0HRuOz2Xo2
XrCvkR/cDDcZqrUKZkyVl/wUxMyE7Rokti5R1zw7gt8q0B4ZMVzm6IbwJAfzNYhL
qNyzr6LLaFW0Jv6fSWhoa567UBcFl9vr1pcSXKA64Mlp/a8q2BICZaxAD/5S0JT/
x9rArVosXsY87UAPOc34FwhDwYEo6qOIjzBy3DLXiroEZbYZtghh2hOZI8zArdMe
5b91wiWHnSBoGzuQtp2Ty7YX0LJf+bdeqEYdP2ayqBsiEjH3AVvqO5qKgEN5vzTu
E3DdfErH4t+v5O855Uvi67OmanPmQyB1vVwAWuWK4fphD6Td9rWu6MFQs9FnWQrB
zJuybeVat5pngYUtNC70A3JMaCFzlsguMt3pjXeGi8VLCpdecaFGuZmq1I9fUw6A
1iNRtnJ1X1yWS0KQm3IBl65y7i0hjkbsFagb+3X1qqLBePw0RL399up6r1dvCk03
wEzkt7ix/1xsjhsO+QqHSnRcB6nEj5ZEKmdJ/3UNTgC2pNVOYKxc4Io6niMlZ0xg
fMaYgrYFhY2PPbJSjKA3qV+Di0VFYx+dD2h6cVITkH8sNlrm/f8bGzmAAIBCM042
5NBZvxp6KrkJ4eM4a6NdZ2A4bbhT90ydGGtN6DcATGPAa+xbtvRGPyI2VJocXd7a
1A3qaHwJsu5q3rHiGyjZF6gdYwOkHG3MfpX/PrTxGs/GTcyX4dpGoEKH0rg7Qg6I
D2AQZ2gGAFSd2FbIHaN5TAwW3vMbPL+GPPOEbgIhi9Jk//p4Ik0XwbHrY00OPeFN
KkOvUijR7PWeJWzaf1p00aHyYvIPo0KHvCG303aO+SHjN+7NUNSxjfYdg17eOWSp
bu4o6H8jTV4vz1MKw2jPpVpYRVWQ+AcYf9GYAouQ18eRBHP8TowWOc/l/ho5d66K
3YVFgaVmmSZ2Fa3+LhmrvVfmXi0bRuZxXoxyb4VEvalVf7z+g+vvwxQ2Gyj2wSm0
rZGABRykM5C+RF3coRhqsXjkra3btNQg3I6ahTuwHlA8QM8R97xm337BhsUKW5hP
WfN5i8slrFatRltka/HSyAt7ZN9zn56Wrv9/yzNRPZof/1AuxDmoQH4NcqAzTE8S
p89A8BGelLAhlM0d94HAfRMpLN1q1yFhLcPJFA1b8JIxCA39PBtrm8S1d8f54y2x
JGDjQ3VSAAeqiHWB0EC6kS30ZDJFSyJwOqol5n8UXIMn8KaSSTDS9grpbBnA/uP4
BedU2JZaBTYYr9j/oMSQES5BsBzZiwMbHsxol4GFGGq1MBOvC6bne6JEIj47HHzf
8rIlWoaVhT93prJpL24YxamNIpotxInOvsfdAsGJFxrj88anrfgKFTDym1mEz9yc
BtN/yuTcBV6ZPMii4klPzUIEbS6sqcNnzk6txIoF2wJguFdAl1yeoYxFfOtQrTfM
Ha10YsiDU7qNyCxudd6B3QBwtdQz0mRcZJ8AfzfBYc0Gyc+piaH05uonlDNzut6D
D3NZyu9s12RLbsPNjyimzPtPfhOY2Oz8I2VAyEVial8FrmnjSNHs2Bmu5lcwprbC
BKjYykgnAxDpn8tO4ijwivNLdhEmrAzucphhO7851xcT6TX8bXU4FJAUBTfmP/G+
i5C+LIG0YXU3WJanAR8LiW6eEgmdcffyIgV4kriFzM2EAIETjnwg3trTUovRdKTk
rYoLEDN/rmK22JX765rrstXMq0UD5UbnK7+mVbZz6B6lNx18J1RKa7ISEL+c/+jj
p6FrmkNu690pKaP4ZiN476r/Pjedt1DBzEDYu+A8X1OhBvL5cWGAiSF25bPbwrIG
tghXxShzlrXNt9+Scxwg68ZTXGtACPXuWUBpQpdC5zXkjiqGQ6GmtR5dgHXRSiV1
YzdnbvmzCU+Wwor3u2MWrUPQdsFGs1SsMAvGV7vYix2AmxRypL0mKsdYIwDzS6Jy
Lpf+M95W5fc8bxHWGhhvun6TqCdWmeGJYIOwPdjUYVlRQEveav8XX3kDNiE13Jrt
DCT+64aqLQCWW1XHPFbTlH21/AGlI/jCqDkhnIdIwIeY+xGqagFif4seNwveirsS
6iMbCcx1el+EF2hzfOAIa2K2YGmOsGfrilF7HTlOH7WY03SNEUFXn+xutwbDGjpB
U3VaLLvponi/u7zu8h1nh/6DrSeYiEuz4uOJD6ACKLwr15fjUMHRYfHIrnYv/358
0CSEngQ7Cd6w9CYK6jDNIFcpSAhYQCkv4PWYdpMbfkI/qu3vb6aeCHcyrqjxrUxG
EpSiHu/VcJsyKEEyXTxxMja02GelAxB+1a4bmVDLiv2KB1gvC/n7PvgU9ZZ+wGV/
y7az7bdGeYVxUO4PnWxmnNZBYis67LGuDiXo/hECW/R683DXBT7KfueT01iDRn6+
2+4har4xMowVDeqJU8eUr495OO5ngt88yfopfxlvmtuUs+l17/Myo84N/5iNeZxz
q5Rp6fevjJwN4/IJLOK1vxm7BWxgyCJHWkWvcaO+Pz74x6sz61sx864ixOk/jmge
raMsmW31hmg1G31XfdiSfYtbVTsoqVRipHWrNN/ZOZPH4jDkAJJQQk/9UwhEXsA4
L95qqn3jMUIUS0dDs2qPnVJpfPoYs172gTb8ZQ4sZjo3NLbB0N6ffg1k3hZEGHj5
dzTAQ6JFb8e73dfYMr8TOH6y2oG+TAUtdvUDQzZZj3cOpzaFKOgswzAf1xe2LlrA
oqOl0iKy/S5MdIPlGIEYycn5+9+M3TYG1VDK52HWA1j1NHSCLX5hvKWVCRiiWAJM
6Ku8TlzmJPedguzfV6i/rhphzsCBrZP5LJwyFAW/psj9fPBcXl1MsBTextA2P4hQ
CHn7I/rjfNhWH6J0wKOlzmBDJSuA/JLxpFYpvoJZDQ1noaoB2jlkO8njqqSPDjSO
bBxniTcrl5r+qC801teQm/5bSv0B0Xyqx3L8b8FQcQu2KhU7vIY1TQwHoxzQ6xKc
Y6SH/8QDHkwZ0ulg34+AAHoSXLAZxmwpTA3G7Rfg4jBUxmLmCa0W5Uoi6kff4KVC
yEuAGKG7LPJe0tpJOQ9OATbQKc7M37XQewPQqTW/IBmcBgmI31xxvcc5vBI2iV95
x25OvKf50Eryn/RslToarnFC9vzDq7brIFVc5oqbZ9O+LSvk5eN/PsiSyeb2jOC7
XaA2DS2CwGQeKW+m9tTfUZOQ7jkTU3s11ZRLH8+BqQpRvHbSmSftc2KP947WCDpw
VGs1wCYH9nlLHTKQxNXI25Vglx4alsaX6rL+M87CU6mBJja7pW/OpLbIbHLxvvh4
DD7Z1OpkhXdfiDVE/3AYdeovHlCcYheogEsXCJUOb3yIh/norVULiOrRoyh/aDDx
0AbyJDBf0aqRoe6W5jB71g16BEhRVgkEGVGZTTYm8YKXF4RJ+XTe1fL7AB/eLRwL
2mmj8fn2BzanVazHSLsE8f4HKHQosLusTkFMUoKmtTDTJba4wohdRHUEh3k2wLrB
mb5r3sY9hsRLLtkFrYmIix6OuMf7S545Yn6YCKcnV3wwrjY0gwME+xNO0PRGqBTN
fKCpyPniJe1hX/4pGmsV2Ov3FeeyRH4UqaX9XApU6fJWvqLROFpB3mTGD0IU2yMc
4yGUOlOgE4izFoUV+oJW1xQFFv0cWP0xb6/yHZE2m02UorpV8X0bGShIsDqAXNHa
N9x9a+pArpq4iZtgPXwZyhSVOYDmtI9nzNfmxhfgkTQFoCOele+bap5CYUYSw+Lk
4pcq2EqmUYCiN2LsA8gUlpMfiYi8ilj6Q0AfpgbkSyokhFO6l0dF4s7pAAA4fG4H
V5xiY5rsViNiYBka8En9WYJM5nLAqRBylR9Gj3eQVKLrwGbSCVKEzH5QvdyXjZ32
dfNrJNHWjkTzTKPksHhZ1QTILh2nuz1crJJTSW5fIoIP/hAMC9FRd5txkRP79jJ4
hq8v2puc8ihr6qW3OdMQZ11z4653zbuTVFpZzJCZ3VE3YNABdR9Zq3kcV5lqHeAf
Rg2NUkeAtSZW3xqwkRRKxSQwMMcTwFSAafGlUGvuaqQ784WyYpv07uNmkH4Aaogc
VXUDfpk84lU8WJxQQ/UF1yQluPrAwuEyzOrDuOkS7yHnkjI42nafP18whgPhBr65
11GW2jEVM5ahDC4STbXhS5/kEtI25BN8Nk7v6TKvx089hEXHscyGfiRuxOk8z1FR
U0a/8vn3WVnBEjsSeKrDsi+k9oYoMBg+KMKEHK2OOQr+Xk2hehkoawTphzeVKCK7
G1t6LJ3PvFt0onq0PuWO/oNU40LHYKQauUzK3ol8uQWk3AKH2ph5H23+QMW7Sg6b
hDQ/sKsZ4m3N8Jxb7rHyKaPeRacQ/xfpaDIV1vp/Scglt8SRtSjiMIlj042l7SXR
5gsv3wXOWQ857GrnKV1G/dogZcGK4DCf7hDWz8/eVH2zqcI5ynwZ594yvtBgneGU
28CofKPpF/+EF/nxHBX3i2nkU+xnRxmSi2iwIjVdcxI7I+QlJKM6aWOkgGBgqYPU
JiSQpsglctsaEWbXqnvnejFRE2Vbn1TgFFR8v5a+pM6Rk9fbixc9WpM5Ss6yrduy
u8/FqnLv1KUWs35eyl7syiFtpj/JxfMFDx/Gd9nE7CTY16BsN2RAhu7WKp/UNLhU
G4miTb7U99uxA9/b70RRGwJuigy1SapPiemq13Ax1R0ty2usINUus7A640opASW4
WnHXofAexZamoV5rQHjE4e4DQNvBrYW2GHmvzhGqjKL4EoNTPu+DCq24FZGtUZ6L
NLKyXkqNO7j3b9zXGtD1sgLceN7h/SEeK4pzfb7cMUazutRlXGhDHsztfNVeILt3
YUFagFbUtSh4P75mMrEW0IpDHur9DCEW7kynLhAp2gVQvXpX+GQtuPCKpM6GENmN
FQ7NB60pqvARwiHooHsuIEEi6RlbbrPyiZvfClmVZ62mUTzgeI5IRdBjcbsu1dp/
mDT9YYoRLnB6u4S98pyLsFUggtEPNmS6UDovqgfq8nh9bYOFGEVi+4apVG/+1dd6
yyvWDp+sIJNkaAnnlM+aGW8EpaY0FHbe+qgUIfJv9M1mMOUboNXDL9znNdWlnXKS
fW5JaiMMTaQ2WMQn3nOXYqOlNp9ngAwrHntyXJGpIHCGzzBRNG74uRf7mLd4foxe
pbjh5A2p080b7qAoKYHOj5Up7ZBSESSRBDHugrptdJeqJ1yj0Tv2UUNBhtzCfUud
GQTrZiSRWNqCi6boGGxId22nUaUM8mSOT1YiMgfZbmC7+FfzW3lKlNQm6b31kx5Y
cqAOmSGgEJs/UZWshKFKlyl8yjzb4abPHpiQuJw5bbGBZHu1De/k2DFb3VRo5vi2
WhG15oaIptnOMrxooDnJjKhhZyMNM+F9VFq/nfRWIqGUOcBLhMvNt3+lJv+7Q45K
ZKEHJyXwqKENxGXG17vwtzPQuSjYCD06yIEUHAssed09z8j+OJJrDIZYRzVS709R
hMP0GHB7n/gBQhL/oCUZLm4vRupMGAk4Rw3Gt9TC1XAomqMpk/wgvcAjpfWZNugJ
+L04Ve2MVvG34tPOsqYGqXU/JcdvYRvMruWPnS7jBtY6wVW6tLbcM9Jbo6ysFXr4
iL4MHgN/7krF0n/n1fw4GQ2J1q90mp9LaSYLjwMEiNEuQkufIlQ4VVV0CHpKOsh0
W1xz6gf1HO+LqEs7yVG6MskIKin284EgoXfkde0AEwILmeumYWvnUIGYW1rLSZu4
3IiIh0RXVQWtTFLoteMR9hFuzoVT8ohWl4yVbOQ09t0lMfekV+Aaj/fZoFOqTUrN
DNelES42PLhWfwIo7SNvjAApqgHZU+LPBY843VG7vwFtSCd0LInDRmqS0Tn16iP+
gz6fA1WdUA6YpbW5V7VKnxfSZuDpO1W74p4m1ewAsTEJyvD8s3SVIjNQ/feogwNu
aAIz7RS5JofT3rxs9kvzLWyj+ky4XpsJ+kH8/ojCmsNQHUJfFlqX3G/9/+Sf3X/f
oyykqOZbZ9lKf0BlL1kl7NXanhd93vFoZZTELboTTsACxjkIQlXGwE6X/llSaI6g
MQieCMjsJWTz9JI0uOtjk8vGX4ggodzyIWdeqWVU+O5nJAZmHd0GPVirzuO0/JRZ
E2ldblgjK46wPJ0wub5SXjPZz0jNl8C6wFlTP2XZDkv/3emQcf0Gdb2HDx7S4WxO
TXOhE6aBl1qrwe/5Z1buPx4wOSBfNGZHIOqh6ZqUWDZMWmFc2aOXc5aszcr7OnrK
utQv/Q3f/0X0HllLQXbaG/zQ2ftbiPmWS4xyOnvJ5CyCi59FOM0XlMdOV591xChX
EmaV+erDMco8TZQlOGIMpYryzpWGSavFD1Bbke4euLjoiXZf2dHdsLYx1tb5udol
rKlqepQOoiyCez3vmqEU4g/q5baackgl6O8i8g3EDkw7MxaE4WVI5qqw6bk2Iwwl
HPsW40+WTC6ayUxcjFY2K9vCAFfySZjlBgsGCKUVcvI47KmXie1HEvm5djWneFbo
DWCYEzwRqagYGB/8bx1jNfr3OCOYe+5a4h2pXek8+0ncm/mtmAUxsIzC7ISDyrwx
OU7eF/C12R65HgJmIK+6fdWQjPPDP9CiAuvHhL++GLqDuR5xGs6rtuO+ZEGdI7Nh
d7YH8HIb+ZgHCAramyQhXD+1AF4rQVoIH170nVN8zkQn52xjfJT0RRXCmZIt9CiR
htJxP2ctC0lSJDiWNyAgT6hOBFQzvjug1BPtVfWS7utuG/dttvtz+Gz7wIHY3bol
eONnEVOJkHBZwYluk8VYKc45uqdWtR9V4s6QfZ/9F3s707Rq0AS1d3Ut+wEyBc8s
vHv6LlO1bnmrkGDyVK8ch+pBO6NW/81vcMAyFoFX8957ECXLlC7IAvVYBehPSl9x
sRlMpU7BYOmolLMuSnLzGOxL8JH7pCgqRB9tbRTlfAQT2y6OtS83UK0XvS6L8MyU
BGkq+bHCzmO4iAvFoo82/V0qxanFIJWzbnv2Z32kwjPA7osUu1OkXCQH5b4BOviK
yTXRcp1NpOGLW+kIvPEorHJoyqk6xauan7zwDo9dB0QkfAAOBhMuFtLhstjegcPb
8jJBjv9466aZ0gJLLEjVoUkYyowarMylttuZ5JfhLQmRuacvVreqA1i0k87l5YyM
FQoKMsJvQvfq4fipJ0B1SIZUS0tYiuHroGXDeHTDtY+g+JOXBdQ0BlLAbD8UpIdR
CLAxR+WXlrD52GN38WFhL9iNQEFePdCmHPzGvk8/eS1bNp5qkFnjpMuymd6v0OL0
GGcwASXKdRwnDW+tEo4ZSNH3jdc01iZwnzgHUph31ZzcY3L3ihsCQk4DS3CtTOMM
CnmhjpWMJuL/chc6pXbFbt8LiEswkDoT4fqPx6cUN8LU2dC81HUD2hHPM8c86zCa
WVRCd9FxJ9npK4bN4JyykFcNR2ydh0o0w3I9RWu4xWkqJY7YLImxVDdKBPHsWYqe
tdcpwS00j8tz2AQUVsdp2tkbZ9pbz/xP7VGOV9BKK5p0luL2mYbBw7LkshSAI1Mo
/Dlqc5rOBLYlniZ/jCQmXmkIjpglavnOWgx3nVsO3rci0BdKkFNvXQnu6GO3YbAO
EqW1DCB5z1F8AkwvDf/huwsoXIbmw9CX2w+P2G9BuWk9aY/i6dCJW4nd4awVaAOS
lNJiWhAxlXP1tW1khGKPjvwqB7KWUJ6JWCM9YogKm3K+f/uykDt3DL/4rB+MQoz4
rEsBbSIC8Bf3xYcoLdqEDH23VlMqxJVJrOY1ND4+d4qh3eLorvYVF8OxO3NuKtbE
8n3R3lmdOfo2hxUT9A85N8bfIPY6S7Q4IOnuJsOtr/H9/EfnG221ddOLVl4+q7h0
ILifbHS5q0vasZVgIN6gpnvSCNPuN98nsGlQ3D20SZAcMCMoKi18t3iiI+Ftu+6l
vIoxZTDwoeIKp1oLW0VAQBvlxwwicPR0jlo4Kjs/Z0CHSWy+81GGXXBF4NzvzlL0
vBpYSWMcjrupZg2SYfSR9rAzxGELQS5x+MKWqrdNiilCAF/9Oa6oY7hPJGtJRgj5
5V828poQ2jFktkMpqpHh48XDaCzi9m1XLqcvcK+hdklVYgeLN4IQD0wPTq2XCo49
obIk0LDuQWaCVBBPTCfxKaZ8ahwHKIad00UIcG/K2Hee2NDfbW3xrZV9rTrMALTw
p7m0UVuOs0XehXGlnXeIRJrci94+t5QQO3L+3bzTYvSjtwtYHuKN0XphrYEWEkxf
2EgolGoKQ0UwoS5Mbwqid7CsIuT09O+pPj3rISd93qqXD3MaEy0cX39NGzPbEijd
4qC5JugE7LBFvGm6/xSySOhBSdI1zIsTvhln1kXCH7pb4Ynw+77luf8x8P5LlhSu
8f6OgzViDcJOVcRaL034Q4Y2a2zpG3OWxqtBiU6MRbjhym8S7KW96qblI0lrWazn
ASOFJo1o0RoEpGxvM/jAsZ747rDBAQ9QmNKEKo8+ZBjMlBsJWrb4S2acbvAJTV7P
bco3vxNxIf9Pe/Rw69nlVzBvZl8WPWE47Ckv3861aELUkytMtJLRN3RxBbbtuLP9
UakEchrHo8htiIu2vByYEcKlfQghMlSzo3tFHHYLVZPMmN1d+YwOt41ZXBRasfXF
pP93kRb6eG/wo6p0jBpRLhEnGns+gKG3GoPQENZNl9NpuB0Y0E5QN77vMWN3Wzw1
OR3xudx3UAbCy2pehKeWkHfbaWFEc+pT8uNtEaMnkeM9XDrpLqcdiAQLUENrOaSY
siBBCawf6DYKY25Q2bxDGUhyph02u7I9rosV68IDdvcbZqPfpQXJFS8D+yooYGDn
t7CUJHx5nyedMtfdcOLfrO8p0jX9gJ0KnloZKx8uGwdyHVNXqv2rgdBIKGfwu+Tc
wqZSkrPgQwyd+jJJgudRoP87VayYztpsyPYP4P0lZQwomp6rCrpQu46BRjWH5afN
vMe1tjcJJTwcwTn+wirVwhDmAaH25O8ClAL2HiZ32wisC40B2rHrMkq/3QfBy+w2
47oiZawOf6sSAsnFEkpaSE55SlAzTCX5phr8mE+jnIKVTxqRr9mij2ALkGsjg7PK
waHCeVl9LOepuNWHm9rD6VsO65mnNg/D3ktwhmh67IGM70nhrNgE3WoAEE9m93tw
iIMytlSqzoobVw7cE0kKTVx75Nd2/g85UeSRX2040JdKNYR6+3/nCFONX4xdsX1f
V0VyDjz+WWFZqNBOs+dfd8Il7WbsAdmiFQ3x2X3VCCswQ4hYSdgn0hkAsMOcMQZW
UK5+NhCryzb9lxKsNp3mLCPxjWrBKVzGEbslmJ5dnL7Z6TFWmHZ2SKBSFQWRB+S3
D6/M0bgsVqtt+TENvwns+MUhaqysipZk6Ie8nsXJNMGWslNEibPLGbUxvRgQnsPU
e+Dqs9AvEiKrSxnPx0mThb34owQ4c8G8NzvByUOUcyOF4JBlVICuTmrWrqEOlAcH
TiVVYDuOz1n4lVPdShRhGpCgBGn7jy6JjwPDe7tbmRB5lsTJhwQT4KQTGg6t9Ztf
0tV3YkGkiouA/mOuuBx4j2Y6VESH3lTbIRhK4uvlQVSsPdtnlQvdMo87M2eb4XFw
Sss4euaAtgLd88DgCkeEZ7+YPuLdyfkH1ItR4+5PwBjDX24xcM6Kx+qc7z5erdfL
JLTSImdrCFYm0qB0lR6TOauJPFgJow/7dMy+GngEkfTC86n5KyRxnp4QImMquZp7
QeKqhn9MjEk88jL3T23WO9KZga8HFTKEf4sog8rVXuuv/yxAgCqHMuYeukdI+Ws+
YSCJIRj0RAohJQzuvIVmvw7DQ/FQ/DqidN3ae2LJXnJHfMRweTUE6aMXFaIIJlOk
vV16Zt9Bfiz6ghuE8xLw1L1CCuTIqhgYuiZ4eHi/dLzpRftqLQVNbALEZMoyCFx1
SQ33xbQlEHiKHyuPVP4S43HOZja6udTArJGe9zTQ/DDIT7pDzBIsELW8NW+dyyjl
aWqWJN5D1ZMHVywLGvRXuGAPg4xBrYKQsw3itrnDLmm6QM1yJDV0NtzKU7+625cz
OTfaqGFClLVKDnPWa/g0k+tHfECDon22+kIIVSlbdl9najv7y0ph+fSEJUFMa0K3
j93QjpWR227DBOA8K98s3AonpPepWEs5Gi3HqW4azfv44GDrXaInn2rO3k3nhB1V
Q0l/vtak+NO9ty/KGByc/YNOQ6+TTefZy9b8nn7kN7PzJSeR9miafCA70l2nnznK
NBNfdIMubZJbZfpZLKXBSiU3cmz0FCL7qOSgpS8O33D5hAuGb4ZESWmsr1PEpGP+
URO4MIRqKoBGpQeZAgDaUkeR4MzVDsvRQf5WqvrBR/ypXZSdsO43VJrmVhGcGEyc
fcONAaSCfgYnI4p10ZgC7oyX3ed2M+fZK87yM+OAd11kkaZQVkFBYQ3eK7J0Fb6v
eBsyeCBkoyLoHHLfMeMax/gJdWPzysiQhrbliEafnk4PdgzkS5G3IVx+jdu1OcHS
q6yXPY/pWWxZldQ3GVAobLw0lyLT8O26masAx8wcJ8XgLEYZlmjgdUnoPUNOX7Vq
1XFgafvz3veL3KEfMvYc60X0Jh6u9IS1mprxP4JTq2VcfA5Jp4acdGseklqcTZm6
tunLGdWv5ZS9a2/4y52Q4yeNzqLVG+lEQN1BUo8RSSDH2/Yo/FjK7tidkqAblRX2
Unug7akbbmGzTmqwwG8NdY3fzcmkYCr1nHLhD76NoTYdo4/R8A8rE0gJRSCwWiau
q3vAo5TbucZ84O5wx+Mr9ROoYCr3Zn1PYuFcGTXsGA8xL/cMMWTgetw9TmvkfF3h
UEh1xdwhUJgxIsLj5IJgLWF0+Lbpp50SmyEvs1ISl/Naap2r51dBDVNCnUfMjzW+
6u3uNknc8aI+uKGs++ff2aoI4RLM20yZD0LBMPSvlm2DMit+7CyjbVNBiDjTKLo7
kXedovvPXkK0uvvVbrE9pa3cIcKKKs/ioXvpeGelQ6XbNj6ZFi7ntfYiniiN5Xqq
SMiCmfG6GdEB1B4JbVP3ADQ9E08xBpO7cgk37PT4lX6RBchwZyDunFv95ruDvTpN
qH3qJJlijstFXCUHFO2twNWOwBTLEfbDnr1n4EK2jhnmrWEecqLu585bDoiKz3lw
T8W8BrulAlO1MYUry3Kp+uOVvb8s5ypDZ/2uQzwfdTjpOZuPfytV9lZV6Gj1mieF
0pkP5r5WaDZJQZIhEe8y7w/MuIQ0UMsUzjHDT8Te87i+TugUWR5V4Qviw0U9pBnh
xZ7uj4xysK/UJUxC0fzf9TrwRolxukJXXGejsswBxFFV//lY0AseVrycraYIflqc
H3yloQ6JGBiw4l8ovYhaiDGKFG1vq+HIWZ3HtApa0di6WopEEVBoGGl5dXm109uT
7x9w3r1Qv/GzkACxV0l8RQ==
`pragma protect end_protected
